# 
#              Synchronous High Density Single Port SRAM Compiler 
# 
#                    UMC 0.13um L130E Fusion(FSG) Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2005 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http:/www.faraday-tech.com
#   
#       Module Name      : SHUD130_128X32X1BM1
#       Words            : 128
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.01  (pf)
#       Data Slew        : 0.016  (ns)
#       CK Slew          : 0.016  (ns)
#       Power Ring Width : 10  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSC0U_D
#       Memaker          : 200701.1.1
#       Date             : 2009/10/23 10:11:39
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SHUD130_128X32X1BM1
CLASS BLOCK ;
FOREIGN SHUD130_128X32X1BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 750.000 BY 124.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 749.000 118.700 750.000 120.900 ;
  LAYER metal3 ;
  RECT 749.000 118.700 750.000 120.900 ;
  LAYER metal2 ;
  RECT 738.660 118.700 750.000 120.900 ;
  LAYER metal1 ;
  RECT 749.000 118.700 750.000 120.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 115.900 750.000 118.100 ;
  LAYER metal3 ;
  RECT 749.000 115.900 750.000 118.100 ;
  LAYER metal2 ;
  RECT 738.660 115.900 750.000 118.100 ;
  LAYER metal1 ;
  RECT 749.000 115.900 750.000 118.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 113.100 750.000 115.300 ;
  LAYER metal3 ;
  RECT 749.000 113.100 750.000 115.300 ;
  LAYER metal2 ;
  RECT 738.660 113.100 750.000 115.300 ;
  LAYER metal1 ;
  RECT 749.000 113.100 750.000 115.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 7.900 750.000 10.100 ;
  LAYER metal3 ;
  RECT 749.000 7.900 750.000 10.100 ;
  LAYER metal2 ;
  RECT 738.660 7.900 750.000 10.100 ;
  LAYER metal1 ;
  RECT 749.000 7.900 750.000 10.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 5.100 750.000 7.300 ;
  LAYER metal3 ;
  RECT 749.000 5.100 750.000 7.300 ;
  LAYER metal2 ;
  RECT 738.660 5.100 750.000 7.300 ;
  LAYER metal1 ;
  RECT 749.000 5.100 750.000 7.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 2.300 750.000 4.500 ;
  LAYER metal3 ;
  RECT 749.000 2.300 750.000 4.500 ;
  LAYER metal2 ;
  RECT 738.660 2.300 750.000 4.500 ;
  LAYER metal1 ;
  RECT 749.000 2.300 750.000 4.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 118.700 1.000 120.900 ;
  LAYER metal3 ;
  RECT 0.000 118.700 1.000 120.900 ;
  LAYER metal2 ;
  RECT 0.000 118.700 11.600 120.900 ;
  LAYER metal1 ;
  RECT 0.000 118.700 1.000 120.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 115.900 1.000 118.100 ;
  LAYER metal3 ;
  RECT 0.000 115.900 1.000 118.100 ;
  LAYER metal2 ;
  RECT 0.000 115.900 11.600 118.100 ;
  LAYER metal1 ;
  RECT 0.000 115.900 1.000 118.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 113.100 1.000 115.300 ;
  LAYER metal3 ;
  RECT 0.000 113.100 1.000 115.300 ;
  LAYER metal2 ;
  RECT 0.000 113.100 11.600 115.300 ;
  LAYER metal1 ;
  RECT 0.000 113.100 1.000 115.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 7.900 1.000 10.100 ;
  LAYER metal3 ;
  RECT 0.000 7.900 1.000 10.100 ;
  LAYER metal2 ;
  RECT 0.000 7.900 11.600 10.100 ;
  LAYER metal1 ;
  RECT 0.000 7.900 1.000 10.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 5.100 1.000 7.300 ;
  LAYER metal3 ;
  RECT 0.000 5.100 1.000 7.300 ;
  LAYER metal2 ;
  RECT 0.000 5.100 11.600 7.300 ;
  LAYER metal1 ;
  RECT 0.000 5.100 1.000 7.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 2.300 1.000 4.500 ;
  LAYER metal3 ;
  RECT 0.000 2.300 1.000 4.500 ;
  LAYER metal2 ;
  RECT 0.000 2.300 11.600 4.500 ;
  LAYER metal1 ;
  RECT 0.000 2.300 1.000 4.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 744.700 123.000 746.900 124.000 ;
  LAYER metal3 ;
  RECT 744.700 123.000 746.900 124.000 ;
  LAYER metal2 ;
  RECT 744.700 112.560 746.900 124.000 ;
  LAYER metal1 ;
  RECT 744.700 123.000 746.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.900 123.000 744.100 124.000 ;
  LAYER metal3 ;
  RECT 741.900 123.000 744.100 124.000 ;
  LAYER metal2 ;
  RECT 741.900 112.560 744.100 124.000 ;
  LAYER metal1 ;
  RECT 741.900 123.000 744.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 739.100 123.000 741.300 124.000 ;
  LAYER metal3 ;
  RECT 739.100 123.000 741.300 124.000 ;
  LAYER metal2 ;
  RECT 739.100 112.560 741.300 124.000 ;
  LAYER metal1 ;
  RECT 739.100 123.000 741.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.900 123.000 10.100 124.000 ;
  LAYER metal3 ;
  RECT 7.900 123.000 10.100 124.000 ;
  LAYER metal2 ;
  RECT 7.900 112.560 10.100 124.000 ;
  LAYER metal1 ;
  RECT 7.900 123.000 10.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 5.100 123.000 7.300 124.000 ;
  LAYER metal3 ;
  RECT 5.100 123.000 7.300 124.000 ;
  LAYER metal2 ;
  RECT 5.100 112.560 7.300 124.000 ;
  LAYER metal1 ;
  RECT 5.100 123.000 7.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 2.300 123.000 4.500 124.000 ;
  LAYER metal3 ;
  RECT 2.300 123.000 4.500 124.000 ;
  LAYER metal2 ;
  RECT 2.300 112.560 4.500 124.000 ;
  LAYER metal1 ;
  RECT 2.300 123.000 4.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 744.700 0.000 746.900 11.600 ;
  LAYER metal3 ;
  RECT 744.700 0.000 746.900 1.000 ;
  LAYER metal2 ;
  RECT 744.700 0.000 746.900 1.000 ;
  LAYER metal1 ;
  RECT 744.700 0.000 746.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.900 0.000 744.100 11.600 ;
  LAYER metal3 ;
  RECT 741.900 0.000 744.100 1.000 ;
  LAYER metal2 ;
  RECT 741.900 0.000 744.100 1.000 ;
  LAYER metal1 ;
  RECT 741.900 0.000 744.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 739.100 0.000 741.300 11.600 ;
  LAYER metal3 ;
  RECT 739.100 0.000 741.300 1.000 ;
  LAYER metal2 ;
  RECT 739.100 0.000 741.300 1.000 ;
  LAYER metal1 ;
  RECT 739.100 0.000 741.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.900 0.000 10.100 11.600 ;
  LAYER metal3 ;
  RECT 7.900 0.000 10.100 1.000 ;
  LAYER metal2 ;
  RECT 7.900 0.000 10.100 1.000 ;
  LAYER metal1 ;
  RECT 7.900 0.000 10.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 5.100 0.000 7.300 11.600 ;
  LAYER metal3 ;
  RECT 5.100 0.000 7.300 1.000 ;
  LAYER metal2 ;
  RECT 5.100 0.000 7.300 1.000 ;
  LAYER metal1 ;
  RECT 5.100 0.000 7.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 2.300 0.000 4.500 11.600 ;
  LAYER metal3 ;
  RECT 2.300 0.000 4.500 1.000 ;
  LAYER metal2 ;
  RECT 2.300 0.000 4.500 1.000 ;
  LAYER metal1 ;
  RECT 2.300 0.000 4.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 89.500 750.000 91.700 ;
  LAYER metal3 ;
  RECT 749.000 89.500 750.000 91.700 ;
  LAYER metal2 ;
  RECT 738.660 89.500 750.000 91.700 ;
  LAYER metal1 ;
  RECT 749.000 89.500 750.000 91.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 83.900 750.000 86.100 ;
  LAYER metal3 ;
  RECT 749.000 83.900 750.000 86.100 ;
  LAYER metal2 ;
  RECT 738.660 83.900 750.000 86.100 ;
  LAYER metal1 ;
  RECT 749.000 83.900 750.000 86.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 78.300 750.000 80.500 ;
  LAYER metal3 ;
  RECT 749.000 78.300 750.000 80.500 ;
  LAYER metal2 ;
  RECT 738.660 78.300 750.000 80.500 ;
  LAYER metal1 ;
  RECT 749.000 78.300 750.000 80.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 33.500 750.000 35.700 ;
  LAYER metal3 ;
  RECT 749.000 33.500 750.000 35.700 ;
  LAYER metal2 ;
  RECT 738.660 33.500 750.000 35.700 ;
  LAYER metal1 ;
  RECT 749.000 33.500 750.000 35.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 27.900 750.000 30.100 ;
  LAYER metal3 ;
  RECT 749.000 27.900 750.000 30.100 ;
  LAYER metal2 ;
  RECT 738.660 27.900 750.000 30.100 ;
  LAYER metal1 ;
  RECT 749.000 27.900 750.000 30.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 22.300 750.000 24.500 ;
  LAYER metal3 ;
  RECT 749.000 22.300 750.000 24.500 ;
  LAYER metal2 ;
  RECT 738.660 22.300 750.000 24.500 ;
  LAYER metal1 ;
  RECT 749.000 22.300 750.000 24.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 89.500 1.000 91.700 ;
  LAYER metal3 ;
  RECT 0.000 89.500 1.000 91.700 ;
  LAYER metal2 ;
  RECT 0.000 89.500 11.600 91.700 ;
  LAYER metal1 ;
  RECT 0.000 89.500 1.000 91.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 83.900 1.000 86.100 ;
  LAYER metal3 ;
  RECT 0.000 83.900 1.000 86.100 ;
  LAYER metal2 ;
  RECT 0.000 83.900 11.600 86.100 ;
  LAYER metal1 ;
  RECT 0.000 83.900 1.000 86.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 78.300 1.000 80.500 ;
  LAYER metal3 ;
  RECT 0.000 78.300 1.000 80.500 ;
  LAYER metal2 ;
  RECT 0.000 78.300 11.600 80.500 ;
  LAYER metal1 ;
  RECT 0.000 78.300 1.000 80.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 33.500 1.000 35.700 ;
  LAYER metal3 ;
  RECT 0.000 33.500 1.000 35.700 ;
  LAYER metal2 ;
  RECT 0.000 33.500 11.600 35.700 ;
  LAYER metal1 ;
  RECT 0.000 33.500 1.000 35.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.900 1.000 30.100 ;
  LAYER metal3 ;
  RECT 0.000 27.900 1.000 30.100 ;
  LAYER metal2 ;
  RECT 0.000 27.900 11.600 30.100 ;
  LAYER metal1 ;
  RECT 0.000 27.900 1.000 30.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 22.300 1.000 24.500 ;
  LAYER metal3 ;
  RECT 0.000 22.300 1.000 24.500 ;
  LAYER metal2 ;
  RECT 0.000 22.300 11.600 24.500 ;
  LAYER metal1 ;
  RECT 0.000 22.300 1.000 24.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 705.500 123.000 707.700 124.000 ;
  LAYER metal3 ;
  RECT 705.500 123.000 707.700 124.000 ;
  LAYER metal2 ;
  RECT 705.500 112.560 707.700 124.000 ;
  LAYER metal1 ;
  RECT 705.500 123.000 707.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 699.900 123.000 702.100 124.000 ;
  LAYER metal3 ;
  RECT 699.900 123.000 702.100 124.000 ;
  LAYER metal2 ;
  RECT 699.900 112.560 702.100 124.000 ;
  LAYER metal1 ;
  RECT 699.900 123.000 702.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 694.300 123.000 696.500 124.000 ;
  LAYER metal3 ;
  RECT 694.300 123.000 696.500 124.000 ;
  LAYER metal2 ;
  RECT 694.300 112.560 696.500 124.000 ;
  LAYER metal1 ;
  RECT 694.300 123.000 696.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 649.500 123.000 651.700 124.000 ;
  LAYER metal3 ;
  RECT 649.500 123.000 651.700 124.000 ;
  LAYER metal2 ;
  RECT 649.500 112.560 651.700 124.000 ;
  LAYER metal1 ;
  RECT 649.500 123.000 651.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 643.900 123.000 646.100 124.000 ;
  LAYER metal3 ;
  RECT 643.900 123.000 646.100 124.000 ;
  LAYER metal2 ;
  RECT 643.900 112.560 646.100 124.000 ;
  LAYER metal1 ;
  RECT 643.900 123.000 646.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 638.300 123.000 640.500 124.000 ;
  LAYER metal3 ;
  RECT 638.300 123.000 640.500 124.000 ;
  LAYER metal2 ;
  RECT 638.300 112.560 640.500 124.000 ;
  LAYER metal1 ;
  RECT 638.300 123.000 640.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 593.500 123.000 595.700 124.000 ;
  LAYER metal3 ;
  RECT 593.500 123.000 595.700 124.000 ;
  LAYER metal2 ;
  RECT 593.500 112.560 595.700 124.000 ;
  LAYER metal1 ;
  RECT 593.500 123.000 595.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 587.900 123.000 590.100 124.000 ;
  LAYER metal3 ;
  RECT 587.900 123.000 590.100 124.000 ;
  LAYER metal2 ;
  RECT 587.900 112.560 590.100 124.000 ;
  LAYER metal1 ;
  RECT 587.900 123.000 590.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 582.300 123.000 584.500 124.000 ;
  LAYER metal3 ;
  RECT 582.300 123.000 584.500 124.000 ;
  LAYER metal2 ;
  RECT 582.300 112.560 584.500 124.000 ;
  LAYER metal1 ;
  RECT 582.300 123.000 584.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.500 123.000 539.700 124.000 ;
  LAYER metal3 ;
  RECT 537.500 123.000 539.700 124.000 ;
  LAYER metal2 ;
  RECT 537.500 112.560 539.700 124.000 ;
  LAYER metal1 ;
  RECT 537.500 123.000 539.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 531.900 123.000 534.100 124.000 ;
  LAYER metal3 ;
  RECT 531.900 123.000 534.100 124.000 ;
  LAYER metal2 ;
  RECT 531.900 112.560 534.100 124.000 ;
  LAYER metal1 ;
  RECT 531.900 123.000 534.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 526.300 123.000 528.500 124.000 ;
  LAYER metal3 ;
  RECT 526.300 123.000 528.500 124.000 ;
  LAYER metal2 ;
  RECT 526.300 112.560 528.500 124.000 ;
  LAYER metal1 ;
  RECT 526.300 123.000 528.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 481.500 123.000 483.700 124.000 ;
  LAYER metal3 ;
  RECT 481.500 123.000 483.700 124.000 ;
  LAYER metal2 ;
  RECT 481.500 112.560 483.700 124.000 ;
  LAYER metal1 ;
  RECT 481.500 123.000 483.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 475.900 123.000 478.100 124.000 ;
  LAYER metal3 ;
  RECT 475.900 123.000 478.100 124.000 ;
  LAYER metal2 ;
  RECT 475.900 112.560 478.100 124.000 ;
  LAYER metal1 ;
  RECT 475.900 123.000 478.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 470.300 123.000 472.500 124.000 ;
  LAYER metal3 ;
  RECT 470.300 123.000 472.500 124.000 ;
  LAYER metal2 ;
  RECT 470.300 112.560 472.500 124.000 ;
  LAYER metal1 ;
  RECT 470.300 123.000 472.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 425.500 123.000 427.700 124.000 ;
  LAYER metal3 ;
  RECT 425.500 123.000 427.700 124.000 ;
  LAYER metal2 ;
  RECT 425.500 112.560 427.700 124.000 ;
  LAYER metal1 ;
  RECT 425.500 123.000 427.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 419.900 123.000 422.100 124.000 ;
  LAYER metal3 ;
  RECT 419.900 123.000 422.100 124.000 ;
  LAYER metal2 ;
  RECT 419.900 112.560 422.100 124.000 ;
  LAYER metal1 ;
  RECT 419.900 123.000 422.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 414.300 123.000 416.500 124.000 ;
  LAYER metal3 ;
  RECT 414.300 123.000 416.500 124.000 ;
  LAYER metal2 ;
  RECT 414.300 112.560 416.500 124.000 ;
  LAYER metal1 ;
  RECT 414.300 123.000 416.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 369.500 123.000 371.700 124.000 ;
  LAYER metal3 ;
  RECT 369.500 123.000 371.700 124.000 ;
  LAYER metal2 ;
  RECT 369.500 112.560 371.700 124.000 ;
  LAYER metal1 ;
  RECT 369.500 123.000 371.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.900 123.000 366.100 124.000 ;
  LAYER metal3 ;
  RECT 363.900 123.000 366.100 124.000 ;
  LAYER metal2 ;
  RECT 363.900 112.560 366.100 124.000 ;
  LAYER metal1 ;
  RECT 363.900 123.000 366.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 358.300 123.000 360.500 124.000 ;
  LAYER metal3 ;
  RECT 358.300 123.000 360.500 124.000 ;
  LAYER metal2 ;
  RECT 358.300 112.560 360.500 124.000 ;
  LAYER metal1 ;
  RECT 358.300 123.000 360.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 313.500 123.000 315.700 124.000 ;
  LAYER metal3 ;
  RECT 313.500 123.000 315.700 124.000 ;
  LAYER metal2 ;
  RECT 313.500 112.560 315.700 124.000 ;
  LAYER metal1 ;
  RECT 313.500 123.000 315.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.900 123.000 310.100 124.000 ;
  LAYER metal3 ;
  RECT 307.900 123.000 310.100 124.000 ;
  LAYER metal2 ;
  RECT 307.900 112.560 310.100 124.000 ;
  LAYER metal1 ;
  RECT 307.900 123.000 310.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.300 123.000 304.500 124.000 ;
  LAYER metal3 ;
  RECT 302.300 123.000 304.500 124.000 ;
  LAYER metal2 ;
  RECT 302.300 112.560 304.500 124.000 ;
  LAYER metal1 ;
  RECT 302.300 123.000 304.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 257.500 123.000 259.700 124.000 ;
  LAYER metal3 ;
  RECT 257.500 123.000 259.700 124.000 ;
  LAYER metal2 ;
  RECT 257.500 112.560 259.700 124.000 ;
  LAYER metal1 ;
  RECT 257.500 123.000 259.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 251.900 123.000 254.100 124.000 ;
  LAYER metal3 ;
  RECT 251.900 123.000 254.100 124.000 ;
  LAYER metal2 ;
  RECT 251.900 112.560 254.100 124.000 ;
  LAYER metal1 ;
  RECT 251.900 123.000 254.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 246.300 123.000 248.500 124.000 ;
  LAYER metal3 ;
  RECT 246.300 123.000 248.500 124.000 ;
  LAYER metal2 ;
  RECT 246.300 112.560 248.500 124.000 ;
  LAYER metal1 ;
  RECT 246.300 123.000 248.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 201.500 123.000 203.700 124.000 ;
  LAYER metal3 ;
  RECT 201.500 123.000 203.700 124.000 ;
  LAYER metal2 ;
  RECT 201.500 112.560 203.700 124.000 ;
  LAYER metal1 ;
  RECT 201.500 123.000 203.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 195.900 123.000 198.100 124.000 ;
  LAYER metal3 ;
  RECT 195.900 123.000 198.100 124.000 ;
  LAYER metal2 ;
  RECT 195.900 112.560 198.100 124.000 ;
  LAYER metal1 ;
  RECT 195.900 123.000 198.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.300 123.000 192.500 124.000 ;
  LAYER metal3 ;
  RECT 190.300 123.000 192.500 124.000 ;
  LAYER metal2 ;
  RECT 190.300 112.560 192.500 124.000 ;
  LAYER metal1 ;
  RECT 190.300 123.000 192.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 145.500 123.000 147.700 124.000 ;
  LAYER metal3 ;
  RECT 145.500 123.000 147.700 124.000 ;
  LAYER metal2 ;
  RECT 145.500 112.560 147.700 124.000 ;
  LAYER metal1 ;
  RECT 145.500 123.000 147.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 123.000 142.100 124.000 ;
  LAYER metal3 ;
  RECT 139.900 123.000 142.100 124.000 ;
  LAYER metal2 ;
  RECT 139.900 112.560 142.100 124.000 ;
  LAYER metal1 ;
  RECT 139.900 123.000 142.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 134.300 123.000 136.500 124.000 ;
  LAYER metal3 ;
  RECT 134.300 123.000 136.500 124.000 ;
  LAYER metal2 ;
  RECT 134.300 112.560 136.500 124.000 ;
  LAYER metal1 ;
  RECT 134.300 123.000 136.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 89.500 123.000 91.700 124.000 ;
  LAYER metal3 ;
  RECT 89.500 123.000 91.700 124.000 ;
  LAYER metal2 ;
  RECT 89.500 112.560 91.700 124.000 ;
  LAYER metal1 ;
  RECT 89.500 123.000 91.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.900 123.000 86.100 124.000 ;
  LAYER metal3 ;
  RECT 83.900 123.000 86.100 124.000 ;
  LAYER metal2 ;
  RECT 83.900 112.560 86.100 124.000 ;
  LAYER metal1 ;
  RECT 83.900 123.000 86.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 78.300 123.000 80.500 124.000 ;
  LAYER metal3 ;
  RECT 78.300 123.000 80.500 124.000 ;
  LAYER metal2 ;
  RECT 78.300 112.560 80.500 124.000 ;
  LAYER metal1 ;
  RECT 78.300 123.000 80.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.500 123.000 35.700 124.000 ;
  LAYER metal3 ;
  RECT 33.500 123.000 35.700 124.000 ;
  LAYER metal2 ;
  RECT 33.500 112.560 35.700 124.000 ;
  LAYER metal1 ;
  RECT 33.500 123.000 35.700 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.900 123.000 30.100 124.000 ;
  LAYER metal3 ;
  RECT 27.900 123.000 30.100 124.000 ;
  LAYER metal2 ;
  RECT 27.900 112.560 30.100 124.000 ;
  LAYER metal1 ;
  RECT 27.900 123.000 30.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 22.300 123.000 24.500 124.000 ;
  LAYER metal3 ;
  RECT 22.300 123.000 24.500 124.000 ;
  LAYER metal2 ;
  RECT 22.300 112.560 24.500 124.000 ;
  LAYER metal1 ;
  RECT 22.300 123.000 24.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 722.700 0.000 724.900 11.600 ;
  LAYER metal3 ;
  RECT 722.700 0.000 724.900 1.000 ;
  LAYER metal2 ;
  RECT 722.700 0.000 724.900 1.000 ;
  LAYER metal1 ;
  RECT 722.700 0.000 724.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 716.300 0.000 718.500 11.600 ;
  LAYER metal3 ;
  RECT 716.300 0.000 718.500 1.000 ;
  LAYER metal2 ;
  RECT 716.300 0.000 718.500 1.000 ;
  LAYER metal1 ;
  RECT 716.300 0.000 718.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.700 0.000 712.900 11.600 ;
  LAYER metal3 ;
  RECT 710.700 0.000 712.900 1.000 ;
  LAYER metal2 ;
  RECT 710.700 0.000 712.900 1.000 ;
  LAYER metal1 ;
  RECT 710.700 0.000 712.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 655.500 0.000 657.700 11.600 ;
  LAYER metal3 ;
  RECT 655.500 0.000 657.700 1.000 ;
  LAYER metal2 ;
  RECT 655.500 0.000 657.700 1.000 ;
  LAYER metal1 ;
  RECT 655.500 0.000 657.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 649.900 0.000 652.100 11.600 ;
  LAYER metal3 ;
  RECT 649.900 0.000 652.100 1.000 ;
  LAYER metal2 ;
  RECT 649.900 0.000 652.100 1.000 ;
  LAYER metal1 ;
  RECT 649.900 0.000 652.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 643.500 0.000 645.700 11.600 ;
  LAYER metal3 ;
  RECT 643.500 0.000 645.700 1.000 ;
  LAYER metal2 ;
  RECT 643.500 0.000 645.700 1.000 ;
  LAYER metal1 ;
  RECT 643.500 0.000 645.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 590.700 0.000 592.900 11.600 ;
  LAYER metal3 ;
  RECT 590.700 0.000 592.900 1.000 ;
  LAYER metal2 ;
  RECT 590.700 0.000 592.900 1.000 ;
  LAYER metal1 ;
  RECT 590.700 0.000 592.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 585.100 0.000 587.300 11.600 ;
  LAYER metal3 ;
  RECT 585.100 0.000 587.300 1.000 ;
  LAYER metal2 ;
  RECT 585.100 0.000 587.300 1.000 ;
  LAYER metal1 ;
  RECT 585.100 0.000 587.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 573.900 0.000 576.100 11.600 ;
  LAYER metal3 ;
  RECT 573.900 0.000 576.100 1.000 ;
  LAYER metal2 ;
  RECT 573.900 0.000 576.100 1.000 ;
  LAYER metal1 ;
  RECT 573.900 0.000 576.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 520.700 0.000 522.900 11.600 ;
  LAYER metal3 ;
  RECT 520.700 0.000 522.900 1.000 ;
  LAYER metal2 ;
  RECT 520.700 0.000 522.900 1.000 ;
  LAYER metal1 ;
  RECT 520.700 0.000 522.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 511.900 0.000 514.100 11.600 ;
  LAYER metal3 ;
  RECT 511.900 0.000 514.100 1.000 ;
  LAYER metal2 ;
  RECT 511.900 0.000 514.100 1.000 ;
  LAYER metal1 ;
  RECT 511.900 0.000 514.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 506.300 0.000 508.500 11.600 ;
  LAYER metal3 ;
  RECT 506.300 0.000 508.500 1.000 ;
  LAYER metal2 ;
  RECT 506.300 0.000 508.500 1.000 ;
  LAYER metal1 ;
  RECT 506.300 0.000 508.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 448.300 0.000 450.500 11.600 ;
  LAYER metal3 ;
  RECT 448.300 0.000 450.500 1.000 ;
  LAYER metal2 ;
  RECT 448.300 0.000 450.500 1.000 ;
  LAYER metal1 ;
  RECT 448.300 0.000 450.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 442.700 0.000 444.900 11.600 ;
  LAYER metal3 ;
  RECT 442.700 0.000 444.900 1.000 ;
  LAYER metal2 ;
  RECT 442.700 0.000 444.900 1.000 ;
  LAYER metal1 ;
  RECT 442.700 0.000 444.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 436.300 0.000 438.500 11.600 ;
  LAYER metal3 ;
  RECT 436.300 0.000 438.500 1.000 ;
  LAYER metal2 ;
  RECT 436.300 0.000 438.500 1.000 ;
  LAYER metal1 ;
  RECT 436.300 0.000 438.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 383.900 0.000 386.100 11.600 ;
  LAYER metal3 ;
  RECT 383.900 0.000 386.100 1.000 ;
  LAYER metal2 ;
  RECT 383.900 0.000 386.100 1.000 ;
  LAYER metal1 ;
  RECT 383.900 0.000 386.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 369.100 0.000 371.300 11.600 ;
  LAYER metal3 ;
  RECT 369.100 0.000 371.300 1.000 ;
  LAYER metal2 ;
  RECT 369.100 0.000 371.300 1.000 ;
  LAYER metal1 ;
  RECT 369.100 0.000 371.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 361.500 0.000 363.700 11.600 ;
  LAYER metal3 ;
  RECT 361.500 0.000 363.700 1.000 ;
  LAYER metal2 ;
  RECT 361.500 0.000 363.700 1.000 ;
  LAYER metal1 ;
  RECT 361.500 0.000 363.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 305.900 0.000 308.100 11.600 ;
  LAYER metal3 ;
  RECT 305.900 0.000 308.100 1.000 ;
  LAYER metal2 ;
  RECT 305.900 0.000 308.100 1.000 ;
  LAYER metal1 ;
  RECT 305.900 0.000 308.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 297.100 0.000 299.300 11.600 ;
  LAYER metal3 ;
  RECT 297.100 0.000 299.300 1.000 ;
  LAYER metal2 ;
  RECT 297.100 0.000 299.300 1.000 ;
  LAYER metal1 ;
  RECT 297.100 0.000 299.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 291.500 0.000 293.700 11.600 ;
  LAYER metal3 ;
  RECT 291.500 0.000 293.700 1.000 ;
  LAYER metal2 ;
  RECT 291.500 0.000 293.700 1.000 ;
  LAYER metal1 ;
  RECT 291.500 0.000 293.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 236.300 0.000 238.500 11.600 ;
  LAYER metal3 ;
  RECT 236.300 0.000 238.500 1.000 ;
  LAYER metal2 ;
  RECT 236.300 0.000 238.500 1.000 ;
  LAYER metal1 ;
  RECT 236.300 0.000 238.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 230.700 0.000 232.900 11.600 ;
  LAYER metal3 ;
  RECT 230.700 0.000 232.900 1.000 ;
  LAYER metal2 ;
  RECT 230.700 0.000 232.900 1.000 ;
  LAYER metal1 ;
  RECT 230.700 0.000 232.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.300 0.000 226.500 11.600 ;
  LAYER metal3 ;
  RECT 224.300 0.000 226.500 1.000 ;
  LAYER metal2 ;
  RECT 224.300 0.000 226.500 1.000 ;
  LAYER metal1 ;
  RECT 224.300 0.000 226.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 171.500 0.000 173.700 11.600 ;
  LAYER metal3 ;
  RECT 171.500 0.000 173.700 1.000 ;
  LAYER metal2 ;
  RECT 171.500 0.000 173.700 1.000 ;
  LAYER metal1 ;
  RECT 171.500 0.000 173.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 163.500 0.000 165.700 11.600 ;
  LAYER metal3 ;
  RECT 163.500 0.000 165.700 1.000 ;
  LAYER metal2 ;
  RECT 163.500 0.000 165.700 1.000 ;
  LAYER metal1 ;
  RECT 163.500 0.000 165.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 157.100 0.000 159.300 11.600 ;
  LAYER metal3 ;
  RECT 157.100 0.000 159.300 1.000 ;
  LAYER metal2 ;
  RECT 157.100 0.000 159.300 1.000 ;
  LAYER metal1 ;
  RECT 157.100 0.000 159.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 104.300 0.000 106.500 11.600 ;
  LAYER metal3 ;
  RECT 104.300 0.000 106.500 1.000 ;
  LAYER metal2 ;
  RECT 104.300 0.000 106.500 1.000 ;
  LAYER metal1 ;
  RECT 104.300 0.000 106.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 97.900 0.000 100.100 11.600 ;
  LAYER metal3 ;
  RECT 97.900 0.000 100.100 1.000 ;
  LAYER metal2 ;
  RECT 97.900 0.000 100.100 1.000 ;
  LAYER metal1 ;
  RECT 97.900 0.000 100.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.300 0.000 94.500 11.600 ;
  LAYER metal3 ;
  RECT 92.300 0.000 94.500 1.000 ;
  LAYER metal2 ;
  RECT 92.300 0.000 94.500 1.000 ;
  LAYER metal1 ;
  RECT 92.300 0.000 94.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 34.300 0.000 36.500 11.600 ;
  LAYER metal3 ;
  RECT 34.300 0.000 36.500 1.000 ;
  LAYER metal2 ;
  RECT 34.300 0.000 36.500 1.000 ;
  LAYER metal1 ;
  RECT 34.300 0.000 36.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 28.700 0.000 30.900 11.600 ;
  LAYER metal3 ;
  RECT 28.700 0.000 30.900 1.000 ;
  LAYER metal2 ;
  RECT 28.700 0.000 30.900 1.000 ;
  LAYER metal1 ;
  RECT 28.700 0.000 30.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 22.300 0.000 24.500 11.600 ;
  LAYER metal3 ;
  RECT 22.300 0.000 24.500 1.000 ;
  LAYER metal2 ;
  RECT 22.300 0.000 24.500 1.000 ;
  LAYER metal1 ;
  RECT 22.300 0.000 24.500 1.000 ;
 END
END VCC
PIN GND
  DIRECTION INPUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 749.000 108.300 750.000 110.500 ;
  LAYER metal3 ;
  RECT 728.380 108.300 750.000 110.500 ;
  LAYER metal2 ;
  RECT 749.000 108.300 750.000 110.500 ;
  LAYER metal1 ;
  RECT 749.000 108.300 750.000 110.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 105.500 750.000 107.700 ;
  LAYER metal3 ;
  RECT 728.380 105.500 750.000 107.700 ;
  LAYER metal2 ;
  RECT 749.000 105.500 750.000 107.700 ;
  LAYER metal1 ;
  RECT 749.000 105.500 750.000 107.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 102.700 750.000 104.900 ;
  LAYER metal3 ;
  RECT 728.380 102.700 750.000 104.900 ;
  LAYER metal2 ;
  RECT 749.000 102.700 750.000 104.900 ;
  LAYER metal1 ;
  RECT 749.000 102.700 750.000 104.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 17.900 750.000 20.100 ;
  LAYER metal3 ;
  RECT 728.380 17.900 750.000 20.100 ;
  LAYER metal2 ;
  RECT 749.000 17.900 750.000 20.100 ;
  LAYER metal1 ;
  RECT 749.000 17.900 750.000 20.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 15.100 750.000 17.300 ;
  LAYER metal3 ;
  RECT 728.380 15.100 750.000 17.300 ;
  LAYER metal2 ;
  RECT 749.000 15.100 750.000 17.300 ;
  LAYER metal1 ;
  RECT 749.000 15.100 750.000 17.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 12.300 750.000 14.500 ;
  LAYER metal3 ;
  RECT 728.380 12.300 750.000 14.500 ;
  LAYER metal2 ;
  RECT 749.000 12.300 750.000 14.500 ;
  LAYER metal1 ;
  RECT 749.000 12.300 750.000 14.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 108.300 1.000 110.500 ;
  LAYER metal3 ;
  RECT 0.000 108.300 21.880 110.500 ;
  LAYER metal2 ;
  RECT 0.000 108.300 1.000 110.500 ;
  LAYER metal1 ;
  RECT 0.000 108.300 1.000 110.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 105.500 1.000 107.700 ;
  LAYER metal3 ;
  RECT 0.000 105.500 21.880 107.700 ;
  LAYER metal2 ;
  RECT 0.000 105.500 1.000 107.700 ;
  LAYER metal1 ;
  RECT 0.000 105.500 1.000 107.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.700 1.000 104.900 ;
  LAYER metal3 ;
  RECT 0.000 102.700 21.880 104.900 ;
  LAYER metal2 ;
  RECT 0.000 102.700 1.000 104.900 ;
  LAYER metal1 ;
  RECT 0.000 102.700 1.000 104.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 17.900 1.000 20.100 ;
  LAYER metal3 ;
  RECT 0.000 17.900 21.880 20.100 ;
  LAYER metal2 ;
  RECT 0.000 17.900 1.000 20.100 ;
  LAYER metal1 ;
  RECT 0.000 17.900 1.000 20.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 15.100 1.000 17.300 ;
  LAYER metal3 ;
  RECT 0.000 15.100 21.880 17.300 ;
  LAYER metal2 ;
  RECT 0.000 15.100 1.000 17.300 ;
  LAYER metal1 ;
  RECT 0.000 15.100 1.000 17.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.300 1.000 14.500 ;
  LAYER metal3 ;
  RECT 0.000 12.300 21.880 14.500 ;
  LAYER metal2 ;
  RECT 0.000 12.300 1.000 14.500 ;
  LAYER metal1 ;
  RECT 0.000 12.300 1.000 14.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 734.700 123.000 736.900 124.000 ;
  LAYER metal3 ;
  RECT 734.700 102.280 736.900 124.000 ;
  LAYER metal2 ;
  RECT 734.700 123.000 736.900 124.000 ;
  LAYER metal1 ;
  RECT 734.700 123.000 736.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 731.900 123.000 734.100 124.000 ;
  LAYER metal3 ;
  RECT 731.900 102.280 734.100 124.000 ;
  LAYER metal2 ;
  RECT 731.900 123.000 734.100 124.000 ;
  LAYER metal1 ;
  RECT 731.900 123.000 734.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 729.100 123.000 731.300 124.000 ;
  LAYER metal3 ;
  RECT 729.100 102.280 731.300 124.000 ;
  LAYER metal2 ;
  RECT 729.100 123.000 731.300 124.000 ;
  LAYER metal1 ;
  RECT 729.100 123.000 731.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 17.900 123.000 20.100 124.000 ;
  LAYER metal3 ;
  RECT 17.900 102.280 20.100 124.000 ;
  LAYER metal2 ;
  RECT 17.900 123.000 20.100 124.000 ;
  LAYER metal1 ;
  RECT 17.900 123.000 20.100 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 15.100 123.000 17.300 124.000 ;
  LAYER metal3 ;
  RECT 15.100 102.280 17.300 124.000 ;
  LAYER metal2 ;
  RECT 15.100 123.000 17.300 124.000 ;
  LAYER metal1 ;
  RECT 15.100 123.000 17.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.300 123.000 14.500 124.000 ;
  LAYER metal3 ;
  RECT 12.300 102.280 14.500 124.000 ;
  LAYER metal2 ;
  RECT 12.300 123.000 14.500 124.000 ;
  LAYER metal1 ;
  RECT 12.300 123.000 14.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 734.700 0.000 736.900 1.000 ;
  LAYER metal3 ;
  RECT 734.700 0.000 736.900 21.880 ;
  LAYER metal2 ;
  RECT 734.700 0.000 736.900 1.000 ;
  LAYER metal1 ;
  RECT 734.700 0.000 736.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 731.900 0.000 734.100 1.000 ;
  LAYER metal3 ;
  RECT 731.900 0.000 734.100 21.880 ;
  LAYER metal2 ;
  RECT 731.900 0.000 734.100 1.000 ;
  LAYER metal1 ;
  RECT 731.900 0.000 734.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 729.100 0.000 731.300 1.000 ;
  LAYER metal3 ;
  RECT 729.100 0.000 731.300 21.880 ;
  LAYER metal2 ;
  RECT 729.100 0.000 731.300 1.000 ;
  LAYER metal1 ;
  RECT 729.100 0.000 731.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 17.900 0.000 20.100 1.000 ;
  LAYER metal3 ;
  RECT 17.900 0.000 20.100 21.880 ;
  LAYER metal2 ;
  RECT 17.900 0.000 20.100 1.000 ;
  LAYER metal1 ;
  RECT 17.900 0.000 20.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 15.100 0.000 17.300 1.000 ;
  LAYER metal3 ;
  RECT 15.100 0.000 17.300 21.880 ;
  LAYER metal2 ;
  RECT 15.100 0.000 17.300 1.000 ;
  LAYER metal1 ;
  RECT 15.100 0.000 17.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.300 0.000 14.500 1.000 ;
  LAYER metal3 ;
  RECT 12.300 0.000 14.500 21.880 ;
  LAYER metal2 ;
  RECT 12.300 0.000 14.500 1.000 ;
  LAYER metal1 ;
  RECT 12.300 0.000 14.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 92.300 750.000 94.500 ;
  LAYER metal3 ;
  RECT 728.380 92.300 750.000 94.500 ;
  LAYER metal2 ;
  RECT 749.000 92.300 750.000 94.500 ;
  LAYER metal1 ;
  RECT 749.000 92.300 750.000 94.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 86.700 750.000 88.900 ;
  LAYER metal3 ;
  RECT 728.380 86.700 750.000 88.900 ;
  LAYER metal2 ;
  RECT 749.000 86.700 750.000 88.900 ;
  LAYER metal1 ;
  RECT 749.000 86.700 750.000 88.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 81.100 750.000 83.300 ;
  LAYER metal3 ;
  RECT 728.380 81.100 750.000 83.300 ;
  LAYER metal2 ;
  RECT 749.000 81.100 750.000 83.300 ;
  LAYER metal1 ;
  RECT 749.000 81.100 750.000 83.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 36.300 750.000 38.500 ;
  LAYER metal3 ;
  RECT 728.380 36.300 750.000 38.500 ;
  LAYER metal2 ;
  RECT 749.000 36.300 750.000 38.500 ;
  LAYER metal1 ;
  RECT 749.000 36.300 750.000 38.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 30.700 750.000 32.900 ;
  LAYER metal3 ;
  RECT 728.380 30.700 750.000 32.900 ;
  LAYER metal2 ;
  RECT 749.000 30.700 750.000 32.900 ;
  LAYER metal1 ;
  RECT 749.000 30.700 750.000 32.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.000 25.100 750.000 27.300 ;
  LAYER metal3 ;
  RECT 728.380 25.100 750.000 27.300 ;
  LAYER metal2 ;
  RECT 749.000 25.100 750.000 27.300 ;
  LAYER metal1 ;
  RECT 749.000 25.100 750.000 27.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 92.300 1.000 94.500 ;
  LAYER metal3 ;
  RECT 0.000 92.300 21.880 94.500 ;
  LAYER metal2 ;
  RECT 0.000 92.300 1.000 94.500 ;
  LAYER metal1 ;
  RECT 0.000 92.300 1.000 94.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.700 1.000 88.900 ;
  LAYER metal3 ;
  RECT 0.000 86.700 21.880 88.900 ;
  LAYER metal2 ;
  RECT 0.000 86.700 1.000 88.900 ;
  LAYER metal1 ;
  RECT 0.000 86.700 1.000 88.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 81.100 1.000 83.300 ;
  LAYER metal3 ;
  RECT 0.000 81.100 21.880 83.300 ;
  LAYER metal2 ;
  RECT 0.000 81.100 1.000 83.300 ;
  LAYER metal1 ;
  RECT 0.000 81.100 1.000 83.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 36.300 1.000 38.500 ;
  LAYER metal3 ;
  RECT 0.000 36.300 21.880 38.500 ;
  LAYER metal2 ;
  RECT 0.000 36.300 1.000 38.500 ;
  LAYER metal1 ;
  RECT 0.000 36.300 1.000 38.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 30.700 1.000 32.900 ;
  LAYER metal3 ;
  RECT 0.000 30.700 21.880 32.900 ;
  LAYER metal2 ;
  RECT 0.000 30.700 1.000 32.900 ;
  LAYER metal1 ;
  RECT 0.000 30.700 1.000 32.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 25.100 1.000 27.300 ;
  LAYER metal3 ;
  RECT 0.000 25.100 21.880 27.300 ;
  LAYER metal2 ;
  RECT 0.000 25.100 1.000 27.300 ;
  LAYER metal1 ;
  RECT 0.000 25.100 1.000 27.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 708.300 123.000 710.500 124.000 ;
  LAYER metal3 ;
  RECT 708.300 102.280 710.500 124.000 ;
  LAYER metal2 ;
  RECT 708.300 123.000 710.500 124.000 ;
  LAYER metal1 ;
  RECT 708.300 123.000 710.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.700 123.000 704.900 124.000 ;
  LAYER metal3 ;
  RECT 702.700 102.280 704.900 124.000 ;
  LAYER metal2 ;
  RECT 702.700 123.000 704.900 124.000 ;
  LAYER metal1 ;
  RECT 702.700 123.000 704.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 697.100 123.000 699.300 124.000 ;
  LAYER metal3 ;
  RECT 697.100 102.280 699.300 124.000 ;
  LAYER metal2 ;
  RECT 697.100 123.000 699.300 124.000 ;
  LAYER metal1 ;
  RECT 697.100 123.000 699.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 652.300 123.000 654.500 124.000 ;
  LAYER metal3 ;
  RECT 652.300 102.280 654.500 124.000 ;
  LAYER metal2 ;
  RECT 652.300 123.000 654.500 124.000 ;
  LAYER metal1 ;
  RECT 652.300 123.000 654.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 646.700 123.000 648.900 124.000 ;
  LAYER metal3 ;
  RECT 646.700 102.280 648.900 124.000 ;
  LAYER metal2 ;
  RECT 646.700 123.000 648.900 124.000 ;
  LAYER metal1 ;
  RECT 646.700 123.000 648.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.100 123.000 643.300 124.000 ;
  LAYER metal3 ;
  RECT 641.100 102.280 643.300 124.000 ;
  LAYER metal2 ;
  RECT 641.100 123.000 643.300 124.000 ;
  LAYER metal1 ;
  RECT 641.100 123.000 643.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 596.300 123.000 598.500 124.000 ;
  LAYER metal3 ;
  RECT 596.300 102.280 598.500 124.000 ;
  LAYER metal2 ;
  RECT 596.300 123.000 598.500 124.000 ;
  LAYER metal1 ;
  RECT 596.300 123.000 598.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 590.700 123.000 592.900 124.000 ;
  LAYER metal3 ;
  RECT 590.700 102.280 592.900 124.000 ;
  LAYER metal2 ;
  RECT 590.700 123.000 592.900 124.000 ;
  LAYER metal1 ;
  RECT 590.700 123.000 592.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 585.100 123.000 587.300 124.000 ;
  LAYER metal3 ;
  RECT 585.100 102.280 587.300 124.000 ;
  LAYER metal2 ;
  RECT 585.100 123.000 587.300 124.000 ;
  LAYER metal1 ;
  RECT 585.100 123.000 587.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 540.300 123.000 542.500 124.000 ;
  LAYER metal3 ;
  RECT 540.300 102.280 542.500 124.000 ;
  LAYER metal2 ;
  RECT 540.300 123.000 542.500 124.000 ;
  LAYER metal1 ;
  RECT 540.300 123.000 542.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 534.700 123.000 536.900 124.000 ;
  LAYER metal3 ;
  RECT 534.700 102.280 536.900 124.000 ;
  LAYER metal2 ;
  RECT 534.700 123.000 536.900 124.000 ;
  LAYER metal1 ;
  RECT 534.700 123.000 536.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 529.100 123.000 531.300 124.000 ;
  LAYER metal3 ;
  RECT 529.100 102.280 531.300 124.000 ;
  LAYER metal2 ;
  RECT 529.100 123.000 531.300 124.000 ;
  LAYER metal1 ;
  RECT 529.100 123.000 531.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 484.300 123.000 486.500 124.000 ;
  LAYER metal3 ;
  RECT 484.300 102.280 486.500 124.000 ;
  LAYER metal2 ;
  RECT 484.300 123.000 486.500 124.000 ;
  LAYER metal1 ;
  RECT 484.300 123.000 486.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 478.700 123.000 480.900 124.000 ;
  LAYER metal3 ;
  RECT 478.700 102.280 480.900 124.000 ;
  LAYER metal2 ;
  RECT 478.700 123.000 480.900 124.000 ;
  LAYER metal1 ;
  RECT 478.700 123.000 480.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 473.100 123.000 475.300 124.000 ;
  LAYER metal3 ;
  RECT 473.100 102.280 475.300 124.000 ;
  LAYER metal2 ;
  RECT 473.100 123.000 475.300 124.000 ;
  LAYER metal1 ;
  RECT 473.100 123.000 475.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 428.300 123.000 430.500 124.000 ;
  LAYER metal3 ;
  RECT 428.300 102.280 430.500 124.000 ;
  LAYER metal2 ;
  RECT 428.300 123.000 430.500 124.000 ;
  LAYER metal1 ;
  RECT 428.300 123.000 430.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 422.700 123.000 424.900 124.000 ;
  LAYER metal3 ;
  RECT 422.700 102.280 424.900 124.000 ;
  LAYER metal2 ;
  RECT 422.700 123.000 424.900 124.000 ;
  LAYER metal1 ;
  RECT 422.700 123.000 424.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 417.100 123.000 419.300 124.000 ;
  LAYER metal3 ;
  RECT 417.100 102.280 419.300 124.000 ;
  LAYER metal2 ;
  RECT 417.100 123.000 419.300 124.000 ;
  LAYER metal1 ;
  RECT 417.100 123.000 419.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.300 123.000 374.500 124.000 ;
  LAYER metal3 ;
  RECT 372.300 102.280 374.500 124.000 ;
  LAYER metal2 ;
  RECT 372.300 123.000 374.500 124.000 ;
  LAYER metal1 ;
  RECT 372.300 123.000 374.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 366.700 123.000 368.900 124.000 ;
  LAYER metal3 ;
  RECT 366.700 102.280 368.900 124.000 ;
  LAYER metal2 ;
  RECT 366.700 123.000 368.900 124.000 ;
  LAYER metal1 ;
  RECT 366.700 123.000 368.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 361.100 123.000 363.300 124.000 ;
  LAYER metal3 ;
  RECT 361.100 102.280 363.300 124.000 ;
  LAYER metal2 ;
  RECT 361.100 123.000 363.300 124.000 ;
  LAYER metal1 ;
  RECT 361.100 123.000 363.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 316.300 123.000 318.500 124.000 ;
  LAYER metal3 ;
  RECT 316.300 102.280 318.500 124.000 ;
  LAYER metal2 ;
  RECT 316.300 123.000 318.500 124.000 ;
  LAYER metal1 ;
  RECT 316.300 123.000 318.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 310.700 123.000 312.900 124.000 ;
  LAYER metal3 ;
  RECT 310.700 102.280 312.900 124.000 ;
  LAYER metal2 ;
  RECT 310.700 123.000 312.900 124.000 ;
  LAYER metal1 ;
  RECT 310.700 123.000 312.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 305.100 123.000 307.300 124.000 ;
  LAYER metal3 ;
  RECT 305.100 102.280 307.300 124.000 ;
  LAYER metal2 ;
  RECT 305.100 123.000 307.300 124.000 ;
  LAYER metal1 ;
  RECT 305.100 123.000 307.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 260.300 123.000 262.500 124.000 ;
  LAYER metal3 ;
  RECT 260.300 102.280 262.500 124.000 ;
  LAYER metal2 ;
  RECT 260.300 123.000 262.500 124.000 ;
  LAYER metal1 ;
  RECT 260.300 123.000 262.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 254.700 123.000 256.900 124.000 ;
  LAYER metal3 ;
  RECT 254.700 102.280 256.900 124.000 ;
  LAYER metal2 ;
  RECT 254.700 123.000 256.900 124.000 ;
  LAYER metal1 ;
  RECT 254.700 123.000 256.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 249.100 123.000 251.300 124.000 ;
  LAYER metal3 ;
  RECT 249.100 102.280 251.300 124.000 ;
  LAYER metal2 ;
  RECT 249.100 123.000 251.300 124.000 ;
  LAYER metal1 ;
  RECT 249.100 123.000 251.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 204.300 123.000 206.500 124.000 ;
  LAYER metal3 ;
  RECT 204.300 102.280 206.500 124.000 ;
  LAYER metal2 ;
  RECT 204.300 123.000 206.500 124.000 ;
  LAYER metal1 ;
  RECT 204.300 123.000 206.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.700 123.000 200.900 124.000 ;
  LAYER metal3 ;
  RECT 198.700 102.280 200.900 124.000 ;
  LAYER metal2 ;
  RECT 198.700 123.000 200.900 124.000 ;
  LAYER metal1 ;
  RECT 198.700 123.000 200.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 193.100 123.000 195.300 124.000 ;
  LAYER metal3 ;
  RECT 193.100 102.280 195.300 124.000 ;
  LAYER metal2 ;
  RECT 193.100 123.000 195.300 124.000 ;
  LAYER metal1 ;
  RECT 193.100 123.000 195.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.300 123.000 150.500 124.000 ;
  LAYER metal3 ;
  RECT 148.300 102.280 150.500 124.000 ;
  LAYER metal2 ;
  RECT 148.300 123.000 150.500 124.000 ;
  LAYER metal1 ;
  RECT 148.300 123.000 150.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.700 123.000 144.900 124.000 ;
  LAYER metal3 ;
  RECT 142.700 102.280 144.900 124.000 ;
  LAYER metal2 ;
  RECT 142.700 123.000 144.900 124.000 ;
  LAYER metal1 ;
  RECT 142.700 123.000 144.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 137.100 123.000 139.300 124.000 ;
  LAYER metal3 ;
  RECT 137.100 102.280 139.300 124.000 ;
  LAYER metal2 ;
  RECT 137.100 123.000 139.300 124.000 ;
  LAYER metal1 ;
  RECT 137.100 123.000 139.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.300 123.000 94.500 124.000 ;
  LAYER metal3 ;
  RECT 92.300 102.280 94.500 124.000 ;
  LAYER metal2 ;
  RECT 92.300 123.000 94.500 124.000 ;
  LAYER metal1 ;
  RECT 92.300 123.000 94.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 86.700 123.000 88.900 124.000 ;
  LAYER metal3 ;
  RECT 86.700 102.280 88.900 124.000 ;
  LAYER metal2 ;
  RECT 86.700 123.000 88.900 124.000 ;
  LAYER metal1 ;
  RECT 86.700 123.000 88.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 81.100 123.000 83.300 124.000 ;
  LAYER metal3 ;
  RECT 81.100 102.280 83.300 124.000 ;
  LAYER metal2 ;
  RECT 81.100 123.000 83.300 124.000 ;
  LAYER metal1 ;
  RECT 81.100 123.000 83.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 36.300 123.000 38.500 124.000 ;
  LAYER metal3 ;
  RECT 36.300 102.280 38.500 124.000 ;
  LAYER metal2 ;
  RECT 36.300 123.000 38.500 124.000 ;
  LAYER metal1 ;
  RECT 36.300 123.000 38.500 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 30.700 123.000 32.900 124.000 ;
  LAYER metal3 ;
  RECT 30.700 102.280 32.900 124.000 ;
  LAYER metal2 ;
  RECT 30.700 123.000 32.900 124.000 ;
  LAYER metal1 ;
  RECT 30.700 123.000 32.900 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.100 123.000 27.300 124.000 ;
  LAYER metal3 ;
  RECT 25.100 102.280 27.300 124.000 ;
  LAYER metal2 ;
  RECT 25.100 123.000 27.300 124.000 ;
  LAYER metal1 ;
  RECT 25.100 123.000 27.300 124.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 725.500 0.000 727.700 1.000 ;
  LAYER metal3 ;
  RECT 725.500 0.000 727.700 21.880 ;
  LAYER metal2 ;
  RECT 725.500 0.000 727.700 1.000 ;
  LAYER metal1 ;
  RECT 725.500 0.000 727.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.100 0.000 721.300 1.000 ;
  LAYER metal3 ;
  RECT 719.100 0.000 721.300 21.880 ;
  LAYER metal2 ;
  RECT 719.100 0.000 721.300 1.000 ;
  LAYER metal1 ;
  RECT 719.100 0.000 721.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 713.500 0.000 715.700 1.000 ;
  LAYER metal3 ;
  RECT 713.500 0.000 715.700 21.880 ;
  LAYER metal2 ;
  RECT 713.500 0.000 715.700 1.000 ;
  LAYER metal1 ;
  RECT 713.500 0.000 715.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.300 0.000 660.500 1.000 ;
  LAYER metal3 ;
  RECT 658.300 0.000 660.500 21.880 ;
  LAYER metal2 ;
  RECT 658.300 0.000 660.500 1.000 ;
  LAYER metal1 ;
  RECT 658.300 0.000 660.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 652.700 0.000 654.900 1.000 ;
  LAYER metal3 ;
  RECT 652.700 0.000 654.900 21.880 ;
  LAYER metal2 ;
  RECT 652.700 0.000 654.900 1.000 ;
  LAYER metal1 ;
  RECT 652.700 0.000 654.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 647.100 0.000 649.300 1.000 ;
  LAYER metal3 ;
  RECT 647.100 0.000 649.300 21.880 ;
  LAYER metal2 ;
  RECT 647.100 0.000 649.300 1.000 ;
  LAYER metal1 ;
  RECT 647.100 0.000 649.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 593.500 0.000 595.700 1.000 ;
  LAYER metal3 ;
  RECT 593.500 0.000 595.700 21.880 ;
  LAYER metal2 ;
  RECT 593.500 0.000 595.700 1.000 ;
  LAYER metal1 ;
  RECT 593.500 0.000 595.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 587.900 0.000 590.100 1.000 ;
  LAYER metal3 ;
  RECT 587.900 0.000 590.100 21.880 ;
  LAYER metal2 ;
  RECT 587.900 0.000 590.100 1.000 ;
  LAYER metal1 ;
  RECT 587.900 0.000 590.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 579.900 0.000 582.100 1.000 ;
  LAYER metal3 ;
  RECT 579.900 0.000 582.100 21.880 ;
  LAYER metal2 ;
  RECT 579.900 0.000 582.100 1.000 ;
  LAYER metal1 ;
  RECT 579.900 0.000 582.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 524.700 0.000 526.900 1.000 ;
  LAYER metal3 ;
  RECT 524.700 0.000 526.900 21.880 ;
  LAYER metal2 ;
  RECT 524.700 0.000 526.900 1.000 ;
  LAYER metal1 ;
  RECT 524.700 0.000 526.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 517.900 0.000 520.100 1.000 ;
  LAYER metal3 ;
  RECT 517.900 0.000 520.100 21.880 ;
  LAYER metal2 ;
  RECT 517.900 0.000 520.100 1.000 ;
  LAYER metal1 ;
  RECT 517.900 0.000 520.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 509.100 0.000 511.300 1.000 ;
  LAYER metal3 ;
  RECT 509.100 0.000 511.300 21.880 ;
  LAYER metal2 ;
  RECT 509.100 0.000 511.300 1.000 ;
  LAYER metal1 ;
  RECT 509.100 0.000 511.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 451.100 0.000 453.300 1.000 ;
  LAYER metal3 ;
  RECT 451.100 0.000 453.300 21.880 ;
  LAYER metal2 ;
  RECT 451.100 0.000 453.300 1.000 ;
  LAYER metal1 ;
  RECT 451.100 0.000 453.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 445.500 0.000 447.700 1.000 ;
  LAYER metal3 ;
  RECT 445.500 0.000 447.700 21.880 ;
  LAYER metal2 ;
  RECT 445.500 0.000 447.700 1.000 ;
  LAYER metal1 ;
  RECT 445.500 0.000 447.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 439.100 0.000 441.300 1.000 ;
  LAYER metal3 ;
  RECT 439.100 0.000 441.300 21.880 ;
  LAYER metal2 ;
  RECT 439.100 0.000 441.300 1.000 ;
  LAYER metal1 ;
  RECT 439.100 0.000 441.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 386.700 0.000 388.900 1.000 ;
  LAYER metal3 ;
  RECT 386.700 0.000 388.900 21.880 ;
  LAYER metal2 ;
  RECT 386.700 0.000 388.900 1.000 ;
  LAYER metal1 ;
  RECT 386.700 0.000 388.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.100 0.000 383.300 1.000 ;
  LAYER metal3 ;
  RECT 381.100 0.000 383.300 21.880 ;
  LAYER metal2 ;
  RECT 381.100 0.000 383.300 1.000 ;
  LAYER metal1 ;
  RECT 381.100 0.000 383.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 364.300 0.000 366.500 1.000 ;
  LAYER metal3 ;
  RECT 364.300 0.000 366.500 21.880 ;
  LAYER metal2 ;
  RECT 364.300 0.000 366.500 1.000 ;
  LAYER metal1 ;
  RECT 364.300 0.000 366.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 308.700 0.000 310.900 1.000 ;
  LAYER metal3 ;
  RECT 308.700 0.000 310.900 21.880 ;
  LAYER metal2 ;
  RECT 308.700 0.000 310.900 1.000 ;
  LAYER metal1 ;
  RECT 308.700 0.000 310.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 299.900 0.000 302.100 1.000 ;
  LAYER metal3 ;
  RECT 299.900 0.000 302.100 21.880 ;
  LAYER metal2 ;
  RECT 299.900 0.000 302.100 1.000 ;
  LAYER metal1 ;
  RECT 299.900 0.000 302.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.300 0.000 296.500 1.000 ;
  LAYER metal3 ;
  RECT 294.300 0.000 296.500 21.880 ;
  LAYER metal2 ;
  RECT 294.300 0.000 296.500 1.000 ;
  LAYER metal1 ;
  RECT 294.300 0.000 296.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.100 0.000 241.300 1.000 ;
  LAYER metal3 ;
  RECT 239.100 0.000 241.300 21.880 ;
  LAYER metal2 ;
  RECT 239.100 0.000 241.300 1.000 ;
  LAYER metal1 ;
  RECT 239.100 0.000 241.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 233.500 0.000 235.700 1.000 ;
  LAYER metal3 ;
  RECT 233.500 0.000 235.700 21.880 ;
  LAYER metal2 ;
  RECT 233.500 0.000 235.700 1.000 ;
  LAYER metal1 ;
  RECT 233.500 0.000 235.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 227.100 0.000 229.300 1.000 ;
  LAYER metal3 ;
  RECT 227.100 0.000 229.300 21.880 ;
  LAYER metal2 ;
  RECT 227.100 0.000 229.300 1.000 ;
  LAYER metal1 ;
  RECT 227.100 0.000 229.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 174.300 0.000 176.500 1.000 ;
  LAYER metal3 ;
  RECT 174.300 0.000 176.500 21.880 ;
  LAYER metal2 ;
  RECT 174.300 0.000 176.500 1.000 ;
  LAYER metal1 ;
  RECT 174.300 0.000 176.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 168.700 0.000 170.900 1.000 ;
  LAYER metal3 ;
  RECT 168.700 0.000 170.900 21.880 ;
  LAYER metal2 ;
  RECT 168.700 0.000 170.900 1.000 ;
  LAYER metal1 ;
  RECT 168.700 0.000 170.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 159.900 0.000 162.100 1.000 ;
  LAYER metal3 ;
  RECT 159.900 0.000 162.100 21.880 ;
  LAYER metal2 ;
  RECT 159.900 0.000 162.100 1.000 ;
  LAYER metal1 ;
  RECT 159.900 0.000 162.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.900 0.000 110.100 1.000 ;
  LAYER metal3 ;
  RECT 107.900 0.000 110.100 21.880 ;
  LAYER metal2 ;
  RECT 107.900 0.000 110.100 1.000 ;
  LAYER metal1 ;
  RECT 107.900 0.000 110.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 101.500 0.000 103.700 1.000 ;
  LAYER metal3 ;
  RECT 101.500 0.000 103.700 21.880 ;
  LAYER metal2 ;
  RECT 101.500 0.000 103.700 1.000 ;
  LAYER metal1 ;
  RECT 101.500 0.000 103.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 95.100 0.000 97.300 1.000 ;
  LAYER metal3 ;
  RECT 95.100 0.000 97.300 21.880 ;
  LAYER metal2 ;
  RECT 95.100 0.000 97.300 1.000 ;
  LAYER metal1 ;
  RECT 95.100 0.000 97.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 37.100 0.000 39.300 1.000 ;
  LAYER metal3 ;
  RECT 37.100 0.000 39.300 21.880 ;
  LAYER metal2 ;
  RECT 37.100 0.000 39.300 1.000 ;
  LAYER metal1 ;
  RECT 37.100 0.000 39.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 31.500 0.000 33.700 1.000 ;
  LAYER metal3 ;
  RECT 31.500 0.000 33.700 21.880 ;
  LAYER metal2 ;
  RECT 31.500 0.000 33.700 1.000 ;
  LAYER metal1 ;
  RECT 31.500 0.000 33.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.900 0.000 28.100 1.000 ;
  LAYER metal3 ;
  RECT 25.900 0.000 28.100 21.880 ;
  LAYER metal2 ;
  RECT 25.900 0.000 28.100 1.000 ;
  LAYER metal1 ;
  RECT 25.900 0.000 28.100 1.000 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 721.600 0.000 722.400 1.000 ;
  LAYER metal3 ;
  RECT 721.600 0.000 722.400 1.000 ;
  LAYER metal2 ;
  RECT 721.600 0.000 722.400 1.000 ;
  LAYER metal1 ;
  RECT 721.600 0.000 722.400 1.000 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 706.800 0.000 707.600 1.000 ;
  LAYER metal3 ;
  RECT 706.800 0.000 707.600 1.000 ;
  LAYER metal2 ;
  RECT 706.800 0.000 707.600 1.000 ;
  LAYER metal1 ;
  RECT 706.800 0.000 707.600 1.000 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 701.600 0.000 702.400 1.000 ;
  LAYER metal3 ;
  RECT 701.600 0.000 702.400 1.000 ;
  LAYER metal2 ;
  RECT 701.600 0.000 702.400 1.000 ;
  LAYER metal1 ;
  RECT 701.600 0.000 702.400 1.000 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 687.200 0.000 688.000 1.000 ;
  LAYER metal3 ;
  RECT 687.200 0.000 688.000 1.000 ;
  LAYER metal2 ;
  RECT 687.200 0.000 688.000 1.000 ;
  LAYER metal1 ;
  RECT 687.200 0.000 688.000 1.000 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 680.800 0.000 681.600 1.000 ;
  LAYER metal3 ;
  RECT 680.800 0.000 681.600 1.000 ;
  LAYER metal2 ;
  RECT 680.800 0.000 681.600 1.000 ;
  LAYER metal1 ;
  RECT 680.800 0.000 681.600 1.000 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER metal3 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER metal2 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER metal1 ;
  RECT 666.000 0.000 666.800 1.000 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 660.800 0.000 661.600 1.000 ;
  LAYER metal3 ;
  RECT 660.800 0.000 661.600 1.000 ;
  LAYER metal2 ;
  RECT 660.800 0.000 661.600 1.000 ;
  LAYER metal1 ;
  RECT 660.800 0.000 661.600 1.000 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 646.000 0.000 646.800 1.000 ;
  LAYER metal3 ;
  RECT 646.000 0.000 646.800 1.000 ;
  LAYER metal2 ;
  RECT 646.000 0.000 646.800 1.000 ;
  LAYER metal1 ;
  RECT 646.000 0.000 646.800 1.000 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 639.600 0.000 640.400 1.000 ;
  LAYER metal3 ;
  RECT 639.600 0.000 640.400 1.000 ;
  LAYER metal2 ;
  RECT 639.600 0.000 640.400 1.000 ;
  LAYER metal1 ;
  RECT 639.600 0.000 640.400 1.000 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 625.200 0.000 626.000 1.000 ;
  LAYER metal3 ;
  RECT 625.200 0.000 626.000 1.000 ;
  LAYER metal2 ;
  RECT 625.200 0.000 626.000 1.000 ;
  LAYER metal1 ;
  RECT 625.200 0.000 626.000 1.000 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 620.000 0.000 620.800 1.000 ;
  LAYER metal3 ;
  RECT 620.000 0.000 620.800 1.000 ;
  LAYER metal2 ;
  RECT 620.000 0.000 620.800 1.000 ;
  LAYER metal1 ;
  RECT 620.000 0.000 620.800 1.000 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 605.200 0.000 606.000 1.000 ;
  LAYER metal3 ;
  RECT 605.200 0.000 606.000 1.000 ;
  LAYER metal2 ;
  RECT 605.200 0.000 606.000 1.000 ;
  LAYER metal1 ;
  RECT 605.200 0.000 606.000 1.000 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 598.800 0.000 599.600 1.000 ;
  LAYER metal3 ;
  RECT 598.800 0.000 599.600 1.000 ;
  LAYER metal2 ;
  RECT 598.800 0.000 599.600 1.000 ;
  LAYER metal1 ;
  RECT 598.800 0.000 599.600 1.000 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 584.000 0.000 584.800 1.000 ;
  LAYER metal3 ;
  RECT 584.000 0.000 584.800 1.000 ;
  LAYER metal2 ;
  RECT 584.000 0.000 584.800 1.000 ;
  LAYER metal1 ;
  RECT 584.000 0.000 584.800 1.000 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 578.800 0.000 579.600 1.000 ;
  LAYER metal3 ;
  RECT 578.800 0.000 579.600 1.000 ;
  LAYER metal2 ;
  RECT 578.800 0.000 579.600 1.000 ;
  LAYER metal1 ;
  RECT 578.800 0.000 579.600 1.000 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 564.400 0.000 565.200 1.000 ;
  LAYER metal3 ;
  RECT 564.400 0.000 565.200 1.000 ;
  LAYER metal2 ;
  RECT 564.400 0.000 565.200 1.000 ;
  LAYER metal1 ;
  RECT 564.400 0.000 565.200 1.000 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 558.000 0.000 558.800 1.000 ;
  LAYER metal3 ;
  RECT 558.000 0.000 558.800 1.000 ;
  LAYER metal2 ;
  RECT 558.000 0.000 558.800 1.000 ;
  LAYER metal1 ;
  RECT 558.000 0.000 558.800 1.000 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 543.200 0.000 544.000 1.000 ;
  LAYER metal3 ;
  RECT 543.200 0.000 544.000 1.000 ;
  LAYER metal2 ;
  RECT 543.200 0.000 544.000 1.000 ;
  LAYER metal1 ;
  RECT 543.200 0.000 544.000 1.000 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 538.000 0.000 538.800 1.000 ;
  LAYER metal3 ;
  RECT 538.000 0.000 538.800 1.000 ;
  LAYER metal2 ;
  RECT 538.000 0.000 538.800 1.000 ;
  LAYER metal1 ;
  RECT 538.000 0.000 538.800 1.000 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 523.600 0.000 524.400 1.000 ;
  LAYER metal3 ;
  RECT 523.600 0.000 524.400 1.000 ;
  LAYER metal2 ;
  RECT 523.600 0.000 524.400 1.000 ;
  LAYER metal1 ;
  RECT 523.600 0.000 524.400 1.000 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 516.800 0.000 517.600 1.000 ;
  LAYER metal3 ;
  RECT 516.800 0.000 517.600 1.000 ;
  LAYER metal2 ;
  RECT 516.800 0.000 517.600 1.000 ;
  LAYER metal1 ;
  RECT 516.800 0.000 517.600 1.000 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 502.400 0.000 503.200 1.000 ;
  LAYER metal3 ;
  RECT 502.400 0.000 503.200 1.000 ;
  LAYER metal2 ;
  RECT 502.400 0.000 503.200 1.000 ;
  LAYER metal1 ;
  RECT 502.400 0.000 503.200 1.000 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 497.200 0.000 498.000 1.000 ;
  LAYER metal3 ;
  RECT 497.200 0.000 498.000 1.000 ;
  LAYER metal2 ;
  RECT 497.200 0.000 498.000 1.000 ;
  LAYER metal1 ;
  RECT 497.200 0.000 498.000 1.000 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 482.400 0.000 483.200 1.000 ;
  LAYER metal3 ;
  RECT 482.400 0.000 483.200 1.000 ;
  LAYER metal2 ;
  RECT 482.400 0.000 483.200 1.000 ;
  LAYER metal1 ;
  RECT 482.400 0.000 483.200 1.000 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 476.000 0.000 476.800 1.000 ;
  LAYER metal3 ;
  RECT 476.000 0.000 476.800 1.000 ;
  LAYER metal2 ;
  RECT 476.000 0.000 476.800 1.000 ;
  LAYER metal1 ;
  RECT 476.000 0.000 476.800 1.000 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 461.600 0.000 462.400 1.000 ;
  LAYER metal3 ;
  RECT 461.600 0.000 462.400 1.000 ;
  LAYER metal2 ;
  RECT 461.600 0.000 462.400 1.000 ;
  LAYER metal1 ;
  RECT 461.600 0.000 462.400 1.000 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 456.000 0.000 456.800 1.000 ;
  LAYER metal3 ;
  RECT 456.000 0.000 456.800 1.000 ;
  LAYER metal2 ;
  RECT 456.000 0.000 456.800 1.000 ;
  LAYER metal1 ;
  RECT 456.000 0.000 456.800 1.000 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 441.600 0.000 442.400 1.000 ;
  LAYER metal3 ;
  RECT 441.600 0.000 442.400 1.000 ;
  LAYER metal2 ;
  RECT 441.600 0.000 442.400 1.000 ;
  LAYER metal1 ;
  RECT 441.600 0.000 442.400 1.000 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 435.200 0.000 436.000 1.000 ;
  LAYER metal3 ;
  RECT 435.200 0.000 436.000 1.000 ;
  LAYER metal2 ;
  RECT 435.200 0.000 436.000 1.000 ;
  LAYER metal1 ;
  RECT 435.200 0.000 436.000 1.000 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 420.400 0.000 421.200 1.000 ;
  LAYER metal3 ;
  RECT 420.400 0.000 421.200 1.000 ;
  LAYER metal2 ;
  RECT 420.400 0.000 421.200 1.000 ;
  LAYER metal1 ;
  RECT 420.400 0.000 421.200 1.000 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 415.200 0.000 416.000 1.000 ;
  LAYER metal3 ;
  RECT 415.200 0.000 416.000 1.000 ;
  LAYER metal2 ;
  RECT 415.200 0.000 416.000 1.000 ;
  LAYER metal1 ;
  RECT 415.200 0.000 416.000 1.000 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 400.800 0.000 401.600 1.000 ;
  LAYER metal3 ;
  RECT 400.800 0.000 401.600 1.000 ;
  LAYER metal2 ;
  RECT 400.800 0.000 401.600 1.000 ;
  LAYER metal1 ;
  RECT 400.800 0.000 401.600 1.000 ;
 END
END DI16
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 380.000 0.000 380.800 1.000 ;
  LAYER metal3 ;
  RECT 380.000 0.000 380.800 1.000 ;
  LAYER metal2 ;
  RECT 380.000 0.000 380.800 1.000 ;
  LAYER metal1 ;
  RECT 380.000 0.000 380.800 1.000 ;
 END
END A3
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 378.800 0.000 379.600 1.000 ;
  LAYER metal3 ;
  RECT 378.800 0.000 379.600 1.000 ;
  LAYER metal2 ;
  RECT 378.800 0.000 379.600 1.000 ;
  LAYER metal1 ;
  RECT 378.800 0.000 379.600 1.000 ;
 END
END A1
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 377.600 0.000 378.400 1.000 ;
  LAYER metal3 ;
  RECT 377.600 0.000 378.400 1.000 ;
  LAYER metal2 ;
  RECT 377.600 0.000 378.400 1.000 ;
  LAYER metal1 ;
  RECT 377.600 0.000 378.400 1.000 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER metal3 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER metal2 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER metal1 ;
  RECT 376.400 0.000 377.200 1.000 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 375.200 0.000 376.000 1.000 ;
  LAYER metal3 ;
  RECT 375.200 0.000 376.000 1.000 ;
  LAYER metal2 ;
  RECT 375.200 0.000 376.000 1.000 ;
  LAYER metal1 ;
  RECT 375.200 0.000 376.000 1.000 ;
 END
END A2
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 374.000 0.000 374.800 1.000 ;
  LAYER metal3 ;
  RECT 374.000 0.000 374.800 1.000 ;
  LAYER metal2 ;
  RECT 374.000 0.000 374.800 1.000 ;
  LAYER metal1 ;
  RECT 374.000 0.000 374.800 1.000 ;
 END
END A0
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.009 ;
 PORT
  LAYER metal4 ;
  RECT 372.000 0.000 372.800 1.000 ;
  LAYER metal3 ;
  RECT 372.000 0.000 372.800 1.000 ;
  LAYER metal2 ;
  RECT 372.000 0.000 372.800 1.000 ;
  LAYER metal1 ;
  RECT 372.000 0.000 372.800 1.000 ;
 END
END WEB
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.036 ;
 PORT
  LAYER metal4 ;
  RECT 368.000 0.000 368.800 1.000 ;
  LAYER metal3 ;
  RECT 368.000 0.000 368.800 1.000 ;
  LAYER metal2 ;
  RECT 368.000 0.000 368.800 1.000 ;
  LAYER metal1 ;
  RECT 368.000 0.000 368.800 1.000 ;
 END
END CK
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 360.400 0.000 361.200 1.000 ;
  LAYER metal3 ;
  RECT 360.400 0.000 361.200 1.000 ;
  LAYER metal2 ;
  RECT 360.400 0.000 361.200 1.000 ;
  LAYER metal1 ;
  RECT 360.400 0.000 361.200 1.000 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 358.000 0.000 358.800 1.000 ;
  LAYER metal3 ;
  RECT 358.000 0.000 358.800 1.000 ;
  LAYER metal2 ;
  RECT 358.000 0.000 358.800 1.000 ;
  LAYER metal1 ;
  RECT 358.000 0.000 358.800 1.000 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.016 ;
 PORT
  LAYER metal4 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER metal3 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER metal2 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER metal1 ;
  RECT 355.200 0.000 356.000 1.000 ;
 END
END A6
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 346.000 0.000 346.800 1.000 ;
  LAYER metal3 ;
  RECT 346.000 0.000 346.800 1.000 ;
  LAYER metal2 ;
  RECT 346.000 0.000 346.800 1.000 ;
  LAYER metal1 ;
  RECT 346.000 0.000 346.800 1.000 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 331.200 0.000 332.000 1.000 ;
  LAYER metal3 ;
  RECT 331.200 0.000 332.000 1.000 ;
  LAYER metal2 ;
  RECT 331.200 0.000 332.000 1.000 ;
  LAYER metal1 ;
  RECT 331.200 0.000 332.000 1.000 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 326.000 0.000 326.800 1.000 ;
  LAYER metal3 ;
  RECT 326.000 0.000 326.800 1.000 ;
  LAYER metal2 ;
  RECT 326.000 0.000 326.800 1.000 ;
  LAYER metal1 ;
  RECT 326.000 0.000 326.800 1.000 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 311.200 0.000 312.000 1.000 ;
  LAYER metal3 ;
  RECT 311.200 0.000 312.000 1.000 ;
  LAYER metal2 ;
  RECT 311.200 0.000 312.000 1.000 ;
  LAYER metal1 ;
  RECT 311.200 0.000 312.000 1.000 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 304.800 0.000 305.600 1.000 ;
  LAYER metal3 ;
  RECT 304.800 0.000 305.600 1.000 ;
  LAYER metal2 ;
  RECT 304.800 0.000 305.600 1.000 ;
  LAYER metal1 ;
  RECT 304.800 0.000 305.600 1.000 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 290.400 0.000 291.200 1.000 ;
  LAYER metal3 ;
  RECT 290.400 0.000 291.200 1.000 ;
  LAYER metal2 ;
  RECT 290.400 0.000 291.200 1.000 ;
  LAYER metal1 ;
  RECT 290.400 0.000 291.200 1.000 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 285.200 0.000 286.000 1.000 ;
  LAYER metal3 ;
  RECT 285.200 0.000 286.000 1.000 ;
  LAYER metal2 ;
  RECT 285.200 0.000 286.000 1.000 ;
  LAYER metal1 ;
  RECT 285.200 0.000 286.000 1.000 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 270.400 0.000 271.200 1.000 ;
  LAYER metal3 ;
  RECT 270.400 0.000 271.200 1.000 ;
  LAYER metal2 ;
  RECT 270.400 0.000 271.200 1.000 ;
  LAYER metal1 ;
  RECT 270.400 0.000 271.200 1.000 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 264.000 0.000 264.800 1.000 ;
  LAYER metal3 ;
  RECT 264.000 0.000 264.800 1.000 ;
  LAYER metal2 ;
  RECT 264.000 0.000 264.800 1.000 ;
  LAYER metal1 ;
  RECT 264.000 0.000 264.800 1.000 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 249.200 0.000 250.000 1.000 ;
  LAYER metal3 ;
  RECT 249.200 0.000 250.000 1.000 ;
  LAYER metal2 ;
  RECT 249.200 0.000 250.000 1.000 ;
  LAYER metal1 ;
  RECT 249.200 0.000 250.000 1.000 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 244.000 0.000 244.800 1.000 ;
  LAYER metal3 ;
  RECT 244.000 0.000 244.800 1.000 ;
  LAYER metal2 ;
  RECT 244.000 0.000 244.800 1.000 ;
  LAYER metal1 ;
  RECT 244.000 0.000 244.800 1.000 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 229.600 0.000 230.400 1.000 ;
  LAYER metal3 ;
  RECT 229.600 0.000 230.400 1.000 ;
  LAYER metal2 ;
  RECT 229.600 0.000 230.400 1.000 ;
  LAYER metal1 ;
  RECT 229.600 0.000 230.400 1.000 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 223.200 0.000 224.000 1.000 ;
  LAYER metal3 ;
  RECT 223.200 0.000 224.000 1.000 ;
  LAYER metal2 ;
  RECT 223.200 0.000 224.000 1.000 ;
  LAYER metal1 ;
  RECT 223.200 0.000 224.000 1.000 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 208.400 0.000 209.200 1.000 ;
  LAYER metal3 ;
  RECT 208.400 0.000 209.200 1.000 ;
  LAYER metal2 ;
  RECT 208.400 0.000 209.200 1.000 ;
  LAYER metal1 ;
  RECT 208.400 0.000 209.200 1.000 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 203.200 0.000 204.000 1.000 ;
  LAYER metal3 ;
  RECT 203.200 0.000 204.000 1.000 ;
  LAYER metal2 ;
  RECT 203.200 0.000 204.000 1.000 ;
  LAYER metal1 ;
  RECT 203.200 0.000 204.000 1.000 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 188.400 0.000 189.200 1.000 ;
  LAYER metal3 ;
  RECT 188.400 0.000 189.200 1.000 ;
  LAYER metal2 ;
  RECT 188.400 0.000 189.200 1.000 ;
  LAYER metal1 ;
  RECT 188.400 0.000 189.200 1.000 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 182.000 0.000 182.800 1.000 ;
  LAYER metal3 ;
  RECT 182.000 0.000 182.800 1.000 ;
  LAYER metal2 ;
  RECT 182.000 0.000 182.800 1.000 ;
  LAYER metal1 ;
  RECT 182.000 0.000 182.800 1.000 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 167.600 0.000 168.400 1.000 ;
  LAYER metal3 ;
  RECT 167.600 0.000 168.400 1.000 ;
  LAYER metal2 ;
  RECT 167.600 0.000 168.400 1.000 ;
  LAYER metal1 ;
  RECT 167.600 0.000 168.400 1.000 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 162.400 0.000 163.200 1.000 ;
  LAYER metal3 ;
  RECT 162.400 0.000 163.200 1.000 ;
  LAYER metal2 ;
  RECT 162.400 0.000 163.200 1.000 ;
  LAYER metal1 ;
  RECT 162.400 0.000 163.200 1.000 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 147.600 0.000 148.400 1.000 ;
  LAYER metal3 ;
  RECT 147.600 0.000 148.400 1.000 ;
  LAYER metal2 ;
  RECT 147.600 0.000 148.400 1.000 ;
  LAYER metal1 ;
  RECT 147.600 0.000 148.400 1.000 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 141.200 0.000 142.000 1.000 ;
  LAYER metal3 ;
  RECT 141.200 0.000 142.000 1.000 ;
  LAYER metal2 ;
  RECT 141.200 0.000 142.000 1.000 ;
  LAYER metal1 ;
  RECT 141.200 0.000 142.000 1.000 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 126.400 0.000 127.200 1.000 ;
  LAYER metal3 ;
  RECT 126.400 0.000 127.200 1.000 ;
  LAYER metal2 ;
  RECT 126.400 0.000 127.200 1.000 ;
  LAYER metal1 ;
  RECT 126.400 0.000 127.200 1.000 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 121.200 0.000 122.000 1.000 ;
  LAYER metal3 ;
  RECT 121.200 0.000 122.000 1.000 ;
  LAYER metal2 ;
  RECT 121.200 0.000 122.000 1.000 ;
  LAYER metal1 ;
  RECT 121.200 0.000 122.000 1.000 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 106.800 0.000 107.600 1.000 ;
  LAYER metal3 ;
  RECT 106.800 0.000 107.600 1.000 ;
  LAYER metal2 ;
  RECT 106.800 0.000 107.600 1.000 ;
  LAYER metal1 ;
  RECT 106.800 0.000 107.600 1.000 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal3 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal2 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal1 ;
  RECT 100.400 0.000 101.200 1.000 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 85.600 0.000 86.400 1.000 ;
  LAYER metal3 ;
  RECT 85.600 0.000 86.400 1.000 ;
  LAYER metal2 ;
  RECT 85.600 0.000 86.400 1.000 ;
  LAYER metal1 ;
  RECT 85.600 0.000 86.400 1.000 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal3 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal2 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal1 ;
  RECT 80.400 0.000 81.200 1.000 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 66.000 0.000 66.800 1.000 ;
  LAYER metal3 ;
  RECT 66.000 0.000 66.800 1.000 ;
  LAYER metal2 ;
  RECT 66.000 0.000 66.800 1.000 ;
  LAYER metal1 ;
  RECT 66.000 0.000 66.800 1.000 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal3 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal2 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal1 ;
  RECT 59.200 0.000 60.000 1.000 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 44.800 0.000 45.600 1.000 ;
  LAYER metal3 ;
  RECT 44.800 0.000 45.600 1.000 ;
  LAYER metal2 ;
  RECT 44.800 0.000 45.600 1.000 ;
  LAYER metal1 ;
  RECT 44.800 0.000 45.600 1.000 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 39.600 0.000 40.400 1.000 ;
  LAYER metal3 ;
  RECT 39.600 0.000 40.400 1.000 ;
  LAYER metal2 ;
  RECT 39.600 0.000 40.400 1.000 ;
  LAYER metal1 ;
  RECT 39.600 0.000 40.400 1.000 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 24.800 0.000 25.600 1.000 ;
  LAYER metal3 ;
  RECT 24.800 0.000 25.600 1.000 ;
  LAYER metal2 ;
  RECT 24.800 0.000 25.600 1.000 ;
  LAYER metal1 ;
  RECT 24.800 0.000 25.600 1.000 ;
 END
END DI0
OBS
  LAYER via4 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER via3 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER via2 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER via ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER metal5 SPACING 0.280 ;
  RECT 20.160 75.940 354.360 104.000 ;
  RECT 392.700 75.940 730.100 104.000 ;
  LAYER metal4 SPACING 0.280 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER metal3 SPACING 0.280 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER metal2 SPACING 0.280 ;
  RECT 0.000 0.200 750.000 124.000 ;
  LAYER metal1 SPACING 0.260 ;
  RECT 0.000 0.200 750.000 124.000 ;
END
END SHUD130_128X32X1BM1
END LIBRARY



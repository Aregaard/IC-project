# 
#              Synchronous Via-1 ROM Compiler 
# 
#                    UMC 0.13um High Speed Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2005 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http:/www.faraday-tech.com
#   
#       Module Name      : SPUD130_512X14BM1A
#       Words            : 512
#       Bits             : 14
#       Aspect Ratio     : 1
#       Output Loading   : 0.01  (pf)
#       Data Slew        : 0.016  (ns)
#       CK Slew          : 0.016  (ns)
#       Power Ring Width : 10  (um)
#       ROM Code File    : /home/piraten/isael/ic-project09/matlab/RomCoeff.txt
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSC0U_D
#       Memaker          : 200701.1.1
#       Date             : 2009/10/23 10:39:18
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SPUD130_512X14BM1A
CLASS BLOCK ;
FOREIGN SPUD130_512X14BM1A 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 230.400 BY 96.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 219.070 90.700 230.400 92.900 ;
  LAYER metal3 ;
  RECT 229.400 90.700 230.400 92.900 ;
  LAYER metal2 ;
  RECT 229.400 90.700 230.400 92.900 ;
  LAYER metal1 ;
  RECT 229.400 90.700 230.400 92.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 87.900 230.400 90.100 ;
  LAYER metal3 ;
  RECT 229.400 87.900 230.400 90.100 ;
  LAYER metal2 ;
  RECT 229.400 87.900 230.400 90.100 ;
  LAYER metal1 ;
  RECT 229.400 87.900 230.400 90.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 85.100 230.400 87.300 ;
  LAYER metal3 ;
  RECT 229.400 85.100 230.400 87.300 ;
  LAYER metal2 ;
  RECT 229.400 85.100 230.400 87.300 ;
  LAYER metal1 ;
  RECT 229.400 85.100 230.400 87.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 7.900 230.400 10.100 ;
  LAYER metal3 ;
  RECT 229.400 7.900 230.400 10.100 ;
  LAYER metal2 ;
  RECT 229.400 7.900 230.400 10.100 ;
  LAYER metal1 ;
  RECT 229.400 7.900 230.400 10.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 5.100 230.400 7.300 ;
  LAYER metal3 ;
  RECT 229.400 5.100 230.400 7.300 ;
  LAYER metal2 ;
  RECT 229.400 5.100 230.400 7.300 ;
  LAYER metal1 ;
  RECT 229.400 5.100 230.400 7.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 2.300 230.400 4.500 ;
  LAYER metal3 ;
  RECT 229.400 2.300 230.400 4.500 ;
  LAYER metal2 ;
  RECT 229.400 2.300 230.400 4.500 ;
  LAYER metal1 ;
  RECT 229.400 2.300 230.400 4.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.700 11.600 92.900 ;
  LAYER metal3 ;
  RECT 0.000 90.700 1.000 92.900 ;
  LAYER metal2 ;
  RECT 0.000 90.700 1.000 92.900 ;
  LAYER metal1 ;
  RECT 0.000 90.700 1.000 92.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 87.900 11.600 90.100 ;
  LAYER metal3 ;
  RECT 0.000 87.900 1.000 90.100 ;
  LAYER metal2 ;
  RECT 0.000 87.900 1.000 90.100 ;
  LAYER metal1 ;
  RECT 0.000 87.900 1.000 90.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 85.100 11.600 87.300 ;
  LAYER metal3 ;
  RECT 0.000 85.100 1.000 87.300 ;
  LAYER metal2 ;
  RECT 0.000 85.100 1.000 87.300 ;
  LAYER metal1 ;
  RECT 0.000 85.100 1.000 87.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 7.900 11.600 10.100 ;
  LAYER metal3 ;
  RECT 0.000 7.900 1.000 10.100 ;
  LAYER metal2 ;
  RECT 0.000 7.900 1.000 10.100 ;
  LAYER metal1 ;
  RECT 0.000 7.900 1.000 10.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 5.100 11.600 7.300 ;
  LAYER metal3 ;
  RECT 0.000 5.100 1.000 7.300 ;
  LAYER metal2 ;
  RECT 0.000 5.100 1.000 7.300 ;
  LAYER metal1 ;
  RECT 0.000 5.100 1.000 7.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 2.300 11.600 4.500 ;
  LAYER metal3 ;
  RECT 0.000 2.300 1.000 4.500 ;
  LAYER metal2 ;
  RECT 0.000 2.300 1.000 4.500 ;
  LAYER metal1 ;
  RECT 0.000 2.300 1.000 4.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 225.100 84.720 227.300 96.000 ;
  LAYER metal3 ;
  RECT 225.100 95.000 227.300 96.000 ;
  LAYER metal2 ;
  RECT 225.100 95.000 227.300 96.000 ;
  LAYER metal1 ;
  RECT 225.100 95.000 227.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.300 84.720 224.500 96.000 ;
  LAYER metal3 ;
  RECT 222.300 95.000 224.500 96.000 ;
  LAYER metal2 ;
  RECT 222.300 95.000 224.500 96.000 ;
  LAYER metal1 ;
  RECT 222.300 95.000 224.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.500 84.720 221.700 96.000 ;
  LAYER metal3 ;
  RECT 219.500 95.000 221.700 96.000 ;
  LAYER metal2 ;
  RECT 219.500 95.000 221.700 96.000 ;
  LAYER metal1 ;
  RECT 219.500 95.000 221.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.900 84.720 10.100 96.000 ;
  LAYER metal3 ;
  RECT 7.900 95.000 10.100 96.000 ;
  LAYER metal2 ;
  RECT 7.900 95.000 10.100 96.000 ;
  LAYER metal1 ;
  RECT 7.900 95.000 10.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 5.100 84.720 7.300 96.000 ;
  LAYER metal3 ;
  RECT 5.100 95.000 7.300 96.000 ;
  LAYER metal2 ;
  RECT 5.100 95.000 7.300 96.000 ;
  LAYER metal1 ;
  RECT 5.100 95.000 7.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 2.300 84.720 4.500 96.000 ;
  LAYER metal3 ;
  RECT 2.300 95.000 4.500 96.000 ;
  LAYER metal2 ;
  RECT 2.300 95.000 4.500 96.000 ;
  LAYER metal1 ;
  RECT 2.300 95.000 4.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 225.100 0.000 227.300 11.600 ;
  LAYER metal3 ;
  RECT 225.100 0.000 227.300 1.000 ;
  LAYER metal2 ;
  RECT 225.100 0.000 227.300 1.000 ;
  LAYER metal1 ;
  RECT 225.100 0.000 227.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.300 0.000 224.500 11.600 ;
  LAYER metal3 ;
  RECT 222.300 0.000 224.500 1.000 ;
  LAYER metal2 ;
  RECT 222.300 0.000 224.500 1.000 ;
  LAYER metal1 ;
  RECT 222.300 0.000 224.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.500 0.000 221.700 11.600 ;
  LAYER metal3 ;
  RECT 219.500 0.000 221.700 1.000 ;
  LAYER metal2 ;
  RECT 219.500 0.000 221.700 1.000 ;
  LAYER metal1 ;
  RECT 219.500 0.000 221.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.900 0.000 10.100 11.600 ;
  LAYER metal3 ;
  RECT 7.900 0.000 10.100 1.000 ;
  LAYER metal2 ;
  RECT 7.900 0.000 10.100 1.000 ;
  LAYER metal1 ;
  RECT 7.900 0.000 10.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 5.100 0.000 7.300 11.600 ;
  LAYER metal3 ;
  RECT 5.100 0.000 7.300 1.000 ;
  LAYER metal2 ;
  RECT 5.100 0.000 7.300 1.000 ;
  LAYER metal1 ;
  RECT 5.100 0.000 7.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 2.300 0.000 4.500 11.600 ;
  LAYER metal3 ;
  RECT 2.300 0.000 4.500 1.000 ;
  LAYER metal2 ;
  RECT 2.300 0.000 4.500 1.000 ;
  LAYER metal1 ;
  RECT 2.300 0.000 4.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 33.500 230.400 35.700 ;
  LAYER metal3 ;
  RECT 229.400 33.500 230.400 35.700 ;
  LAYER metal2 ;
  RECT 229.400 33.500 230.400 35.700 ;
  LAYER metal1 ;
  RECT 229.400 33.500 230.400 35.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 27.900 230.400 30.100 ;
  LAYER metal3 ;
  RECT 229.400 27.900 230.400 30.100 ;
  LAYER metal2 ;
  RECT 229.400 27.900 230.400 30.100 ;
  LAYER metal1 ;
  RECT 229.400 27.900 230.400 30.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 219.070 22.300 230.400 24.500 ;
  LAYER metal3 ;
  RECT 229.400 22.300 230.400 24.500 ;
  LAYER metal2 ;
  RECT 229.400 22.300 230.400 24.500 ;
  LAYER metal1 ;
  RECT 229.400 22.300 230.400 24.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 33.500 11.600 35.700 ;
  LAYER metal3 ;
  RECT 0.000 33.500 1.000 35.700 ;
  LAYER metal2 ;
  RECT 0.000 33.500 1.000 35.700 ;
  LAYER metal1 ;
  RECT 0.000 33.500 1.000 35.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.900 11.600 30.100 ;
  LAYER metal3 ;
  RECT 0.000 27.900 1.000 30.100 ;
  LAYER metal2 ;
  RECT 0.000 27.900 1.000 30.100 ;
  LAYER metal1 ;
  RECT 0.000 27.900 1.000 30.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 22.300 11.600 24.500 ;
  LAYER metal3 ;
  RECT 0.000 22.300 1.000 24.500 ;
  LAYER metal2 ;
  RECT 0.000 22.300 1.000 24.500 ;
  LAYER metal1 ;
  RECT 0.000 22.300 1.000 24.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 201.500 84.720 203.700 96.000 ;
  LAYER metal3 ;
  RECT 201.500 95.000 203.700 96.000 ;
  LAYER metal2 ;
  RECT 201.500 95.000 203.700 96.000 ;
  LAYER metal1 ;
  RECT 201.500 95.000 203.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 195.900 84.720 198.100 96.000 ;
  LAYER metal3 ;
  RECT 195.900 95.000 198.100 96.000 ;
  LAYER metal2 ;
  RECT 195.900 95.000 198.100 96.000 ;
  LAYER metal1 ;
  RECT 195.900 95.000 198.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.300 84.720 192.500 96.000 ;
  LAYER metal3 ;
  RECT 190.300 95.000 192.500 96.000 ;
  LAYER metal2 ;
  RECT 190.300 95.000 192.500 96.000 ;
  LAYER metal1 ;
  RECT 190.300 95.000 192.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 145.500 84.720 147.700 96.000 ;
  LAYER metal3 ;
  RECT 145.500 95.000 147.700 96.000 ;
  LAYER metal2 ;
  RECT 145.500 95.000 147.700 96.000 ;
  LAYER metal1 ;
  RECT 145.500 95.000 147.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 84.720 142.100 96.000 ;
  LAYER metal3 ;
  RECT 139.900 95.000 142.100 96.000 ;
  LAYER metal2 ;
  RECT 139.900 95.000 142.100 96.000 ;
  LAYER metal1 ;
  RECT 139.900 95.000 142.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 134.300 84.720 136.500 96.000 ;
  LAYER metal3 ;
  RECT 134.300 95.000 136.500 96.000 ;
  LAYER metal2 ;
  RECT 134.300 95.000 136.500 96.000 ;
  LAYER metal1 ;
  RECT 134.300 95.000 136.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 89.500 84.720 91.700 96.000 ;
  LAYER metal3 ;
  RECT 89.500 95.000 91.700 96.000 ;
  LAYER metal2 ;
  RECT 89.500 95.000 91.700 96.000 ;
  LAYER metal1 ;
  RECT 89.500 95.000 91.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.900 84.720 86.100 96.000 ;
  LAYER metal3 ;
  RECT 83.900 95.000 86.100 96.000 ;
  LAYER metal2 ;
  RECT 83.900 95.000 86.100 96.000 ;
  LAYER metal1 ;
  RECT 83.900 95.000 86.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 78.300 84.720 80.500 96.000 ;
  LAYER metal3 ;
  RECT 78.300 95.000 80.500 96.000 ;
  LAYER metal2 ;
  RECT 78.300 95.000 80.500 96.000 ;
  LAYER metal1 ;
  RECT 78.300 95.000 80.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.500 84.720 35.700 96.000 ;
  LAYER metal3 ;
  RECT 33.500 95.000 35.700 96.000 ;
  LAYER metal2 ;
  RECT 33.500 95.000 35.700 96.000 ;
  LAYER metal1 ;
  RECT 33.500 95.000 35.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.900 84.720 30.100 96.000 ;
  LAYER metal3 ;
  RECT 27.900 95.000 30.100 96.000 ;
  LAYER metal2 ;
  RECT 27.900 95.000 30.100 96.000 ;
  LAYER metal1 ;
  RECT 27.900 95.000 30.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 22.300 84.720 24.500 96.000 ;
  LAYER metal3 ;
  RECT 22.300 95.000 24.500 96.000 ;
  LAYER metal2 ;
  RECT 22.300 95.000 24.500 96.000 ;
  LAYER metal1 ;
  RECT 22.300 95.000 24.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.100 0.000 205.300 11.600 ;
  LAYER metal3 ;
  RECT 203.100 0.000 205.300 1.000 ;
  LAYER metal2 ;
  RECT 203.100 0.000 205.300 1.000 ;
  LAYER metal1 ;
  RECT 203.100 0.000 205.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 195.500 0.000 197.700 11.600 ;
  LAYER metal3 ;
  RECT 195.500 0.000 197.700 1.000 ;
  LAYER metal2 ;
  RECT 195.500 0.000 197.700 1.000 ;
  LAYER metal1 ;
  RECT 195.500 0.000 197.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 187.900 0.000 190.100 11.600 ;
  LAYER metal3 ;
  RECT 187.900 0.000 190.100 1.000 ;
  LAYER metal2 ;
  RECT 187.900 0.000 190.100 1.000 ;
  LAYER metal1 ;
  RECT 187.900 0.000 190.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.500 0.000 127.700 11.600 ;
  LAYER metal3 ;
  RECT 125.500 0.000 127.700 1.000 ;
  LAYER metal2 ;
  RECT 125.500 0.000 127.700 1.000 ;
  LAYER metal1 ;
  RECT 125.500 0.000 127.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 119.900 0.000 122.100 11.600 ;
  LAYER metal3 ;
  RECT 119.900 0.000 122.100 1.000 ;
  LAYER metal2 ;
  RECT 119.900 0.000 122.100 1.000 ;
  LAYER metal1 ;
  RECT 119.900 0.000 122.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 105.100 0.000 107.300 11.600 ;
  LAYER metal3 ;
  RECT 105.100 0.000 107.300 1.000 ;
  LAYER metal2 ;
  RECT 105.100 0.000 107.300 1.000 ;
  LAYER metal1 ;
  RECT 105.100 0.000 107.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 36.700 0.000 38.900 11.600 ;
  LAYER metal3 ;
  RECT 36.700 0.000 38.900 1.000 ;
  LAYER metal2 ;
  RECT 36.700 0.000 38.900 1.000 ;
  LAYER metal1 ;
  RECT 36.700 0.000 38.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.100 0.000 31.300 11.600 ;
  LAYER metal3 ;
  RECT 29.100 0.000 31.300 1.000 ;
  LAYER metal2 ;
  RECT 29.100 0.000 31.300 1.000 ;
  LAYER metal1 ;
  RECT 29.100 0.000 31.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 22.300 0.000 24.500 11.600 ;
  LAYER metal3 ;
  RECT 22.300 0.000 24.500 1.000 ;
  LAYER metal2 ;
  RECT 22.300 0.000 24.500 1.000 ;
  LAYER metal1 ;
  RECT 22.300 0.000 24.500 1.000 ;
 END
END VCC
PIN GND
  DIRECTION INPUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 229.400 80.700 230.400 82.900 ;
  LAYER metal3 ;
  RECT 208.790 80.700 230.400 82.900 ;
  LAYER metal2 ;
  RECT 229.400 80.700 230.400 82.900 ;
  LAYER metal1 ;
  RECT 229.400 80.700 230.400 82.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 77.900 230.400 80.100 ;
  LAYER metal3 ;
  RECT 208.790 77.900 230.400 80.100 ;
  LAYER metal2 ;
  RECT 229.400 77.900 230.400 80.100 ;
  LAYER metal1 ;
  RECT 229.400 77.900 230.400 80.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 75.100 230.400 77.300 ;
  LAYER metal3 ;
  RECT 208.790 75.100 230.400 77.300 ;
  LAYER metal2 ;
  RECT 229.400 75.100 230.400 77.300 ;
  LAYER metal1 ;
  RECT 229.400 75.100 230.400 77.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 17.900 230.400 20.100 ;
  LAYER metal3 ;
  RECT 208.790 17.900 230.400 20.100 ;
  LAYER metal2 ;
  RECT 229.400 17.900 230.400 20.100 ;
  LAYER metal1 ;
  RECT 229.400 17.900 230.400 20.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 15.100 230.400 17.300 ;
  LAYER metal3 ;
  RECT 208.790 15.100 230.400 17.300 ;
  LAYER metal2 ;
  RECT 229.400 15.100 230.400 17.300 ;
  LAYER metal1 ;
  RECT 229.400 15.100 230.400 17.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 12.300 230.400 14.500 ;
  LAYER metal3 ;
  RECT 208.790 12.300 230.400 14.500 ;
  LAYER metal2 ;
  RECT 229.400 12.300 230.400 14.500 ;
  LAYER metal1 ;
  RECT 229.400 12.300 230.400 14.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 80.700 1.000 82.900 ;
  LAYER metal3 ;
  RECT 0.000 80.700 21.880 82.900 ;
  LAYER metal2 ;
  RECT 0.000 80.700 1.000 82.900 ;
  LAYER metal1 ;
  RECT 0.000 80.700 1.000 82.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 77.900 1.000 80.100 ;
  LAYER metal3 ;
  RECT 0.000 77.900 21.880 80.100 ;
  LAYER metal2 ;
  RECT 0.000 77.900 1.000 80.100 ;
  LAYER metal1 ;
  RECT 0.000 77.900 1.000 80.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 75.100 1.000 77.300 ;
  LAYER metal3 ;
  RECT 0.000 75.100 21.880 77.300 ;
  LAYER metal2 ;
  RECT 0.000 75.100 1.000 77.300 ;
  LAYER metal1 ;
  RECT 0.000 75.100 1.000 77.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 17.900 1.000 20.100 ;
  LAYER metal3 ;
  RECT 0.000 17.900 21.880 20.100 ;
  LAYER metal2 ;
  RECT 0.000 17.900 1.000 20.100 ;
  LAYER metal1 ;
  RECT 0.000 17.900 1.000 20.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 15.100 1.000 17.300 ;
  LAYER metal3 ;
  RECT 0.000 15.100 21.880 17.300 ;
  LAYER metal2 ;
  RECT 0.000 15.100 1.000 17.300 ;
  LAYER metal1 ;
  RECT 0.000 15.100 1.000 17.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.300 1.000 14.500 ;
  LAYER metal3 ;
  RECT 0.000 12.300 21.880 14.500 ;
  LAYER metal2 ;
  RECT 0.000 12.300 1.000 14.500 ;
  LAYER metal1 ;
  RECT 0.000 12.300 1.000 14.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 215.100 95.000 217.300 96.000 ;
  LAYER metal3 ;
  RECT 215.100 74.440 217.300 96.000 ;
  LAYER metal2 ;
  RECT 215.100 95.000 217.300 96.000 ;
  LAYER metal1 ;
  RECT 215.100 95.000 217.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 212.300 95.000 214.500 96.000 ;
  LAYER metal3 ;
  RECT 212.300 74.440 214.500 96.000 ;
  LAYER metal2 ;
  RECT 212.300 95.000 214.500 96.000 ;
  LAYER metal1 ;
  RECT 212.300 95.000 214.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 209.500 95.000 211.700 96.000 ;
  LAYER metal3 ;
  RECT 209.500 74.440 211.700 96.000 ;
  LAYER metal2 ;
  RECT 209.500 95.000 211.700 96.000 ;
  LAYER metal1 ;
  RECT 209.500 95.000 211.700 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 17.900 95.000 20.100 96.000 ;
  LAYER metal3 ;
  RECT 17.900 74.440 20.100 96.000 ;
  LAYER metal2 ;
  RECT 17.900 95.000 20.100 96.000 ;
  LAYER metal1 ;
  RECT 17.900 95.000 20.100 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 15.100 95.000 17.300 96.000 ;
  LAYER metal3 ;
  RECT 15.100 74.440 17.300 96.000 ;
  LAYER metal2 ;
  RECT 15.100 95.000 17.300 96.000 ;
  LAYER metal1 ;
  RECT 15.100 95.000 17.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.300 95.000 14.500 96.000 ;
  LAYER metal3 ;
  RECT 12.300 74.440 14.500 96.000 ;
  LAYER metal2 ;
  RECT 12.300 95.000 14.500 96.000 ;
  LAYER metal1 ;
  RECT 12.300 95.000 14.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 215.100 0.000 217.300 1.000 ;
  LAYER metal3 ;
  RECT 215.100 0.000 217.300 21.880 ;
  LAYER metal2 ;
  RECT 215.100 0.000 217.300 1.000 ;
  LAYER metal1 ;
  RECT 215.100 0.000 217.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 212.300 0.000 214.500 1.000 ;
  LAYER metal3 ;
  RECT 212.300 0.000 214.500 21.880 ;
  LAYER metal2 ;
  RECT 212.300 0.000 214.500 1.000 ;
  LAYER metal1 ;
  RECT 212.300 0.000 214.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 209.500 0.000 211.700 1.000 ;
  LAYER metal3 ;
  RECT 209.500 0.000 211.700 21.880 ;
  LAYER metal2 ;
  RECT 209.500 0.000 211.700 1.000 ;
  LAYER metal1 ;
  RECT 209.500 0.000 211.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 17.900 0.000 20.100 1.000 ;
  LAYER metal3 ;
  RECT 17.900 0.000 20.100 21.880 ;
  LAYER metal2 ;
  RECT 17.900 0.000 20.100 1.000 ;
  LAYER metal1 ;
  RECT 17.900 0.000 20.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 15.100 0.000 17.300 1.000 ;
  LAYER metal3 ;
  RECT 15.100 0.000 17.300 21.880 ;
  LAYER metal2 ;
  RECT 15.100 0.000 17.300 1.000 ;
  LAYER metal1 ;
  RECT 15.100 0.000 17.300 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.300 0.000 14.500 1.000 ;
  LAYER metal3 ;
  RECT 12.300 0.000 14.500 21.880 ;
  LAYER metal2 ;
  RECT 12.300 0.000 14.500 1.000 ;
  LAYER metal1 ;
  RECT 12.300 0.000 14.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 36.300 230.400 38.500 ;
  LAYER metal3 ;
  RECT 208.790 36.300 230.400 38.500 ;
  LAYER metal2 ;
  RECT 229.400 36.300 230.400 38.500 ;
  LAYER metal1 ;
  RECT 229.400 36.300 230.400 38.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 30.700 230.400 32.900 ;
  LAYER metal3 ;
  RECT 208.790 30.700 230.400 32.900 ;
  LAYER metal2 ;
  RECT 229.400 30.700 230.400 32.900 ;
  LAYER metal1 ;
  RECT 229.400 30.700 230.400 32.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.400 25.100 230.400 27.300 ;
  LAYER metal3 ;
  RECT 208.790 25.100 230.400 27.300 ;
  LAYER metal2 ;
  RECT 229.400 25.100 230.400 27.300 ;
  LAYER metal1 ;
  RECT 229.400 25.100 230.400 27.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 36.300 1.000 38.500 ;
  LAYER metal3 ;
  RECT 0.000 36.300 21.880 38.500 ;
  LAYER metal2 ;
  RECT 0.000 36.300 1.000 38.500 ;
  LAYER metal1 ;
  RECT 0.000 36.300 1.000 38.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 30.700 1.000 32.900 ;
  LAYER metal3 ;
  RECT 0.000 30.700 21.880 32.900 ;
  LAYER metal2 ;
  RECT 0.000 30.700 1.000 32.900 ;
  LAYER metal1 ;
  RECT 0.000 30.700 1.000 32.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 25.100 1.000 27.300 ;
  LAYER metal3 ;
  RECT 0.000 25.100 21.880 27.300 ;
  LAYER metal2 ;
  RECT 0.000 25.100 1.000 27.300 ;
  LAYER metal1 ;
  RECT 0.000 25.100 1.000 27.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 204.300 95.000 206.500 96.000 ;
  LAYER metal3 ;
  RECT 204.300 74.440 206.500 96.000 ;
  LAYER metal2 ;
  RECT 204.300 95.000 206.500 96.000 ;
  LAYER metal1 ;
  RECT 204.300 95.000 206.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.700 95.000 200.900 96.000 ;
  LAYER metal3 ;
  RECT 198.700 74.440 200.900 96.000 ;
  LAYER metal2 ;
  RECT 198.700 95.000 200.900 96.000 ;
  LAYER metal1 ;
  RECT 198.700 95.000 200.900 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 193.100 95.000 195.300 96.000 ;
  LAYER metal3 ;
  RECT 193.100 74.440 195.300 96.000 ;
  LAYER metal2 ;
  RECT 193.100 95.000 195.300 96.000 ;
  LAYER metal1 ;
  RECT 193.100 95.000 195.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.300 95.000 150.500 96.000 ;
  LAYER metal3 ;
  RECT 148.300 74.440 150.500 96.000 ;
  LAYER metal2 ;
  RECT 148.300 95.000 150.500 96.000 ;
  LAYER metal1 ;
  RECT 148.300 95.000 150.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.700 95.000 144.900 96.000 ;
  LAYER metal3 ;
  RECT 142.700 74.440 144.900 96.000 ;
  LAYER metal2 ;
  RECT 142.700 95.000 144.900 96.000 ;
  LAYER metal1 ;
  RECT 142.700 95.000 144.900 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 137.100 95.000 139.300 96.000 ;
  LAYER metal3 ;
  RECT 137.100 74.440 139.300 96.000 ;
  LAYER metal2 ;
  RECT 137.100 95.000 139.300 96.000 ;
  LAYER metal1 ;
  RECT 137.100 95.000 139.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.300 95.000 94.500 96.000 ;
  LAYER metal3 ;
  RECT 92.300 74.440 94.500 96.000 ;
  LAYER metal2 ;
  RECT 92.300 95.000 94.500 96.000 ;
  LAYER metal1 ;
  RECT 92.300 95.000 94.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 86.700 95.000 88.900 96.000 ;
  LAYER metal3 ;
  RECT 86.700 74.440 88.900 96.000 ;
  LAYER metal2 ;
  RECT 86.700 95.000 88.900 96.000 ;
  LAYER metal1 ;
  RECT 86.700 95.000 88.900 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 81.100 95.000 83.300 96.000 ;
  LAYER metal3 ;
  RECT 81.100 74.440 83.300 96.000 ;
  LAYER metal2 ;
  RECT 81.100 95.000 83.300 96.000 ;
  LAYER metal1 ;
  RECT 81.100 95.000 83.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 36.300 95.000 38.500 96.000 ;
  LAYER metal3 ;
  RECT 36.300 74.440 38.500 96.000 ;
  LAYER metal2 ;
  RECT 36.300 95.000 38.500 96.000 ;
  LAYER metal1 ;
  RECT 36.300 95.000 38.500 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 30.700 95.000 32.900 96.000 ;
  LAYER metal3 ;
  RECT 30.700 74.440 32.900 96.000 ;
  LAYER metal2 ;
  RECT 30.700 95.000 32.900 96.000 ;
  LAYER metal1 ;
  RECT 30.700 95.000 32.900 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.100 95.000 27.300 96.000 ;
  LAYER metal3 ;
  RECT 25.100 74.440 27.300 96.000 ;
  LAYER metal2 ;
  RECT 25.100 95.000 27.300 96.000 ;
  LAYER metal1 ;
  RECT 25.100 95.000 27.300 96.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 205.900 0.000 208.100 1.000 ;
  LAYER metal3 ;
  RECT 205.900 0.000 208.100 21.880 ;
  LAYER metal2 ;
  RECT 205.900 0.000 208.100 1.000 ;
  LAYER metal1 ;
  RECT 205.900 0.000 208.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.300 0.000 200.500 1.000 ;
  LAYER metal3 ;
  RECT 198.300 0.000 200.500 21.880 ;
  LAYER metal2 ;
  RECT 198.300 0.000 200.500 1.000 ;
  LAYER metal1 ;
  RECT 198.300 0.000 200.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.700 0.000 192.900 1.000 ;
  LAYER metal3 ;
  RECT 190.700 0.000 192.900 21.880 ;
  LAYER metal2 ;
  RECT 190.700 0.000 192.900 1.000 ;
  LAYER metal1 ;
  RECT 190.700 0.000 192.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 130.300 0.000 132.500 1.000 ;
  LAYER metal3 ;
  RECT 130.300 0.000 132.500 21.880 ;
  LAYER metal2 ;
  RECT 130.300 0.000 132.500 1.000 ;
  LAYER metal1 ;
  RECT 130.300 0.000 132.500 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 122.700 0.000 124.900 1.000 ;
  LAYER metal3 ;
  RECT 122.700 0.000 124.900 21.880 ;
  LAYER metal2 ;
  RECT 122.700 0.000 124.900 1.000 ;
  LAYER metal1 ;
  RECT 122.700 0.000 124.900 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.900 0.000 110.100 1.000 ;
  LAYER metal3 ;
  RECT 107.900 0.000 110.100 21.880 ;
  LAYER metal2 ;
  RECT 107.900 0.000 110.100 1.000 ;
  LAYER metal1 ;
  RECT 107.900 0.000 110.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 39.500 0.000 41.700 1.000 ;
  LAYER metal3 ;
  RECT 39.500 0.000 41.700 21.880 ;
  LAYER metal2 ;
  RECT 39.500 0.000 41.700 1.000 ;
  LAYER metal1 ;
  RECT 39.500 0.000 41.700 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 31.900 0.000 34.100 1.000 ;
  LAYER metal3 ;
  RECT 31.900 0.000 34.100 21.880 ;
  LAYER metal2 ;
  RECT 31.900 0.000 34.100 1.000 ;
  LAYER metal1 ;
  RECT 31.900 0.000 34.100 1.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.100 0.000 27.300 1.000 ;
  LAYER metal3 ;
  RECT 25.100 0.000 27.300 21.880 ;
  LAYER metal2 ;
  RECT 25.100 0.000 27.300 1.000 ;
  LAYER metal1 ;
  RECT 25.100 0.000 27.300 1.000 ;
 END
END GND
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 202.000 0.000 202.800 1.000 ;
  LAYER metal3 ;
  RECT 202.000 0.000 202.800 1.000 ;
  LAYER metal2 ;
  RECT 202.000 0.000 202.800 1.000 ;
  LAYER metal1 ;
  RECT 202.000 0.000 202.800 1.000 ;
 END
END DO13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 194.400 0.000 195.200 1.000 ;
  LAYER metal3 ;
  RECT 194.400 0.000 195.200 1.000 ;
  LAYER metal2 ;
  RECT 194.400 0.000 195.200 1.000 ;
  LAYER metal1 ;
  RECT 194.400 0.000 195.200 1.000 ;
 END
END DO12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 186.800 0.000 187.600 1.000 ;
  LAYER metal3 ;
  RECT 186.800 0.000 187.600 1.000 ;
  LAYER metal2 ;
  RECT 186.800 0.000 187.600 1.000 ;
  LAYER metal1 ;
  RECT 186.800 0.000 187.600 1.000 ;
 END
END DO11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 178.400 0.000 179.200 1.000 ;
  LAYER metal3 ;
  RECT 178.400 0.000 179.200 1.000 ;
  LAYER metal2 ;
  RECT 178.400 0.000 179.200 1.000 ;
  LAYER metal1 ;
  RECT 178.400 0.000 179.200 1.000 ;
 END
END DO10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 170.800 0.000 171.600 1.000 ;
  LAYER metal3 ;
  RECT 170.800 0.000 171.600 1.000 ;
  LAYER metal2 ;
  RECT 170.800 0.000 171.600 1.000 ;
  LAYER metal1 ;
  RECT 170.800 0.000 171.600 1.000 ;
 END
END DO9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 162.800 0.000 163.600 1.000 ;
  LAYER metal3 ;
  RECT 162.800 0.000 163.600 1.000 ;
  LAYER metal2 ;
  RECT 162.800 0.000 163.600 1.000 ;
  LAYER metal1 ;
  RECT 162.800 0.000 163.600 1.000 ;
 END
END DO8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 155.200 0.000 156.000 1.000 ;
  LAYER metal3 ;
  RECT 155.200 0.000 156.000 1.000 ;
  LAYER metal2 ;
  RECT 155.200 0.000 156.000 1.000 ;
  LAYER metal1 ;
  RECT 155.200 0.000 156.000 1.000 ;
 END
END DO7
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 138.000 0.000 138.800 1.000 ;
  LAYER metal3 ;
  RECT 138.000 0.000 138.800 1.000 ;
  LAYER metal2 ;
  RECT 138.000 0.000 138.800 1.000 ;
  LAYER metal1 ;
  RECT 138.000 0.000 138.800 1.000 ;
 END
END OE
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 129.200 0.000 130.000 1.000 ;
  LAYER metal3 ;
  RECT 129.200 0.000 130.000 1.000 ;
  LAYER metal2 ;
  RECT 129.200 0.000 130.000 1.000 ;
  LAYER metal1 ;
  RECT 129.200 0.000 130.000 1.000 ;
 END
END CK
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 118.800 0.000 119.600 1.000 ;
  LAYER metal3 ;
  RECT 118.800 0.000 119.600 1.000 ;
  LAYER metal2 ;
  RECT 118.800 0.000 119.600 1.000 ;
  LAYER metal1 ;
  RECT 118.800 0.000 119.600 1.000 ;
 END
END A3
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 115.600 0.000 116.400 1.000 ;
  LAYER metal3 ;
  RECT 115.600 0.000 116.400 1.000 ;
  LAYER metal2 ;
  RECT 115.600 0.000 116.400 1.000 ;
  LAYER metal1 ;
  RECT 115.600 0.000 116.400 1.000 ;
 END
END A2
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.035 ;
 PORT
  LAYER metal4 ;
  RECT 114.000 0.000 114.800 1.000 ;
  LAYER metal3 ;
  RECT 114.000 0.000 114.800 1.000 ;
  LAYER metal2 ;
  RECT 114.000 0.000 114.800 1.000 ;
  LAYER metal1 ;
  RECT 114.000 0.000 114.800 1.000 ;
 END
END CS
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 112.000 0.000 112.800 1.000 ;
  LAYER metal3 ;
  RECT 112.000 0.000 112.800 1.000 ;
  LAYER metal2 ;
  RECT 112.000 0.000 112.800 1.000 ;
  LAYER metal1 ;
  RECT 112.000 0.000 112.800 1.000 ;
 END
END A1
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 104.000 0.000 104.800 1.000 ;
  LAYER metal3 ;
  RECT 104.000 0.000 104.800 1.000 ;
  LAYER metal2 ;
  RECT 104.000 0.000 104.800 1.000 ;
  LAYER metal1 ;
  RECT 104.000 0.000 104.800 1.000 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal3 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal2 ;
  RECT 100.400 0.000 101.200 1.000 ;
  LAYER metal1 ;
  RECT 100.400 0.000 101.200 1.000 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 94.800 0.000 95.600 1.000 ;
  LAYER metal3 ;
  RECT 94.800 0.000 95.600 1.000 ;
  LAYER metal2 ;
  RECT 94.800 0.000 95.600 1.000 ;
  LAYER metal1 ;
  RECT 94.800 0.000 95.600 1.000 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 87.200 0.000 88.000 1.000 ;
  LAYER metal3 ;
  RECT 87.200 0.000 88.000 1.000 ;
  LAYER metal2 ;
  RECT 87.200 0.000 88.000 1.000 ;
  LAYER metal1 ;
  RECT 87.200 0.000 88.000 1.000 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 86.000 0.000 86.800 1.000 ;
  LAYER metal3 ;
  RECT 86.000 0.000 86.800 1.000 ;
  LAYER metal2 ;
  RECT 86.000 0.000 86.800 1.000 ;
  LAYER metal1 ;
  RECT 86.000 0.000 86.800 1.000 ;
 END
END A8
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.015 ;
 PORT
  LAYER metal4 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal3 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal2 ;
  RECT 80.400 0.000 81.200 1.000 ;
  LAYER metal1 ;
  RECT 80.400 0.000 81.200 1.000 ;
 END
END A0
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 74.800 0.000 75.600 1.000 ;
  LAYER metal3 ;
  RECT 74.800 0.000 75.600 1.000 ;
  LAYER metal2 ;
  RECT 74.800 0.000 75.600 1.000 ;
  LAYER metal1 ;
  RECT 74.800 0.000 75.600 1.000 ;
 END
END DO6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 66.800 0.000 67.600 1.000 ;
  LAYER metal3 ;
  RECT 66.800 0.000 67.600 1.000 ;
  LAYER metal2 ;
  RECT 66.800 0.000 67.600 1.000 ;
  LAYER metal1 ;
  RECT 66.800 0.000 67.600 1.000 ;
 END
END DO5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal3 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal2 ;
  RECT 59.200 0.000 60.000 1.000 ;
  LAYER metal1 ;
  RECT 59.200 0.000 60.000 1.000 ;
 END
END DO4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 50.800 0.000 51.600 1.000 ;
  LAYER metal3 ;
  RECT 50.800 0.000 51.600 1.000 ;
  LAYER metal2 ;
  RECT 50.800 0.000 51.600 1.000 ;
  LAYER metal1 ;
  RECT 50.800 0.000 51.600 1.000 ;
 END
END DO3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 43.200 0.000 44.000 1.000 ;
  LAYER metal3 ;
  RECT 43.200 0.000 44.000 1.000 ;
  LAYER metal2 ;
  RECT 43.200 0.000 44.000 1.000 ;
  LAYER metal1 ;
  RECT 43.200 0.000 44.000 1.000 ;
 END
END DO2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 35.600 0.000 36.400 1.000 ;
  LAYER metal3 ;
  RECT 35.600 0.000 36.400 1.000 ;
  LAYER metal2 ;
  RECT 35.600 0.000 36.400 1.000 ;
  LAYER metal1 ;
  RECT 35.600 0.000 36.400 1.000 ;
 END
END DO1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.019 ;
 PORT
  LAYER metal4 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER metal3 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER metal2 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER metal1 ;
  RECT 28.000 0.000 28.800 1.000 ;
 END
END DO0
OBS
  LAYER via3 ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER via2 ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER via ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER metal4 SPACING 0.280 ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER metal3 SPACING 0.280 ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER metal2 SPACING 0.280 ;
  RECT 0.000 0.200 230.400 96.000 ;
  LAYER metal1 SPACING 0.260 ;
  RECT 0.000 0.200 230.400 96.000 ;
END
END SPUD130_512X14BM1A
END LIBRARY


